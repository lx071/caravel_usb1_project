// This is the unpowered netlist.
module usb_top (app_clk,
    reg_ack,
    reg_cs,
    reg_wr,
    usb_clk,
    usb_in_dn,
    usb_in_dp,
    usb_intr_o,
    usb_out_dn,
    usb_out_dp,
    usb_out_tx_oen,
    usb_rstn,
    wbd_clk_int,
    wbd_clk_usb,
    cfg_cska_usb,
    reg_addr,
    reg_be,
    reg_rdata,
    reg_wdata);
 input app_clk;
 output reg_ack;
 input reg_cs;
 input reg_wr;
 input usb_clk;
 input usb_in_dn;
 input usb_in_dp;
 output usb_intr_o;
 output usb_out_dn;
 output usb_out_dp;
 output usb_out_tx_oen;
 input usb_rstn;
 input wbd_clk_int;
 output wbd_clk_usb;
 input [3:0] cfg_cska_usb;
 input [8:0] reg_addr;
 input [3:0] reg_be;
 output [31:0] reg_rdata;
 input [31:0] reg_wdata;

 wire clknet_0_app_clk;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_0_u_usb_host.u_core._171_ ;
 wire \clknet_0_u_usb_host.u_core._172_ ;
 wire \clknet_0_u_usb_host.u_core._178_ ;
 wire \clknet_0_u_usb_host.u_core._183_ ;
 wire \clknet_0_u_usb_host.u_core._184_ ;
 wire \clknet_0_u_usb_host.u_core._185_ ;
 wire \clknet_0_u_usb_host.u_core._186_ ;
 wire \clknet_0_u_usb_host.u_core._192_ ;
 wire \clknet_0_u_usb_host.u_core._193_ ;
 wire \clknet_0_u_usb_host.u_core._200_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0784_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0785_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0786_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_rx._0787_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0721_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0722_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0723_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0724_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0725_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0726_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0727_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0728_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0729_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0730_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0731_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0732_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0733_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0734_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0735_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0736_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0737_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0738_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0739_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0740_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0741_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0742_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0743_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0744_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0745_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0746_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0747_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0748_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0749_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0750_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0751_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0752_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0753_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0754_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0755_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0756_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0757_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0758_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0759_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0760_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0761_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0762_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0763_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0764_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0765_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0766_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0767_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0768_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0769_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0770_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0771_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0772_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0773_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0774_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0775_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0776_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0777_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0778_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0779_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0780_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0781_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0782_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0783_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0784_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0785_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0786_ ;
 wire \clknet_0_u_usb_host.u_core.u_fifo_tx._0787_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._294_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._295_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._296_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._305_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._306_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._307_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._308_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._310_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._311_ ;
 wire \clknet_0_u_usb_host.u_core.u_sie._312_ ;
 wire \clknet_0_u_usb_host.u_phy._173_ ;
 wire \clknet_0_u_usb_host.u_phy._176_ ;
 wire \clknet_0_u_usb_host.u_phy._178_ ;
 wire \clknet_0_u_usb_host.u_phy._179_ ;
 wire \clknet_0_u_usb_host.u_phy._182_ ;
 wire clknet_0_usb_clk;
 wire clknet_1_0__leaf_app_clk;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._171_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._172_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._178_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._183_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._184_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._185_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._186_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._192_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core._193_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._294_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._307_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._308_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._311_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._173_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._176_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._178_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._179_ ;
 wire \clknet_1_0__leaf_u_usb_host.u_phy._182_ ;
 wire clknet_1_1__leaf_app_clk;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._171_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._172_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._178_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._183_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._184_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._185_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._186_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._192_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core._193_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._294_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._307_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._308_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._311_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._173_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._176_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._178_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._179_ ;
 wire \clknet_1_1__leaf_u_usb_host.u_phy._182_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_core._200_ ;
 wire \clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ;
 wire clknet_3_0_0_usb_clk;
 wire clknet_3_1_0_usb_clk;
 wire clknet_3_2_0_usb_clk;
 wire clknet_3_3_0_usb_clk;
 wire clknet_3_4_0_usb_clk;
 wire clknet_3_5_0_usb_clk;
 wire clknet_3_6_0_usb_clk;
 wire clknet_3_7_0_usb_clk;
 wire clknet_leaf_0_usb_clk;
 wire clknet_leaf_10_usb_clk;
 wire clknet_leaf_11_usb_clk;
 wire clknet_leaf_12_usb_clk;
 wire clknet_leaf_13_usb_clk;
 wire clknet_leaf_14_usb_clk;
 wire clknet_leaf_15_usb_clk;
 wire clknet_leaf_16_usb_clk;
 wire clknet_leaf_17_usb_clk;
 wire clknet_leaf_18_usb_clk;
 wire clknet_leaf_19_usb_clk;
 wire clknet_leaf_1_usb_clk;
 wire clknet_leaf_20_usb_clk;
 wire clknet_leaf_21_usb_clk;
 wire clknet_leaf_22_usb_clk;
 wire clknet_leaf_23_usb_clk;
 wire clknet_leaf_24_usb_clk;
 wire clknet_leaf_25_usb_clk;
 wire clknet_leaf_26_usb_clk;
 wire clknet_leaf_27_usb_clk;
 wire clknet_leaf_28_usb_clk;
 wire clknet_leaf_29_usb_clk;
 wire clknet_leaf_2_usb_clk;
 wire clknet_leaf_30_usb_clk;
 wire clknet_leaf_31_usb_clk;
 wire clknet_leaf_32_usb_clk;
 wire clknet_leaf_34_usb_clk;
 wire clknet_leaf_35_usb_clk;
 wire clknet_leaf_36_usb_clk;
 wire clknet_leaf_37_usb_clk;
 wire clknet_leaf_38_usb_clk;
 wire clknet_leaf_39_usb_clk;
 wire clknet_leaf_3_usb_clk;
 wire clknet_leaf_40_usb_clk;
 wire clknet_leaf_42_usb_clk;
 wire clknet_leaf_43_usb_clk;
 wire clknet_leaf_44_usb_clk;
 wire clknet_leaf_45_usb_clk;
 wire clknet_leaf_46_usb_clk;
 wire clknet_leaf_47_usb_clk;
 wire clknet_leaf_49_usb_clk;
 wire clknet_leaf_4_usb_clk;
 wire clknet_leaf_51_usb_clk;
 wire clknet_leaf_53_usb_clk;
 wire clknet_leaf_54_usb_clk;
 wire clknet_leaf_55_usb_clk;
 wire clknet_leaf_56_usb_clk;
 wire clknet_leaf_57_usb_clk;
 wire clknet_leaf_58_usb_clk;
 wire clknet_leaf_59_usb_clk;
 wire clknet_leaf_5_usb_clk;
 wire clknet_leaf_6_usb_clk;
 wire clknet_leaf_7_usb_clk;
 wire clknet_leaf_8_usb_clk;
 wire clknet_leaf_9_usb_clk;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net17;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net18;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net19;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net2;
 wire net20;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net21;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net22;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net23;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \u_skew_usb.clk_d1 ;
 wire \u_skew_usb.clk_d10 ;
 wire \u_skew_usb.clk_d11 ;
 wire \u_skew_usb.clk_d12 ;
 wire \u_skew_usb.clk_d13 ;
 wire \u_skew_usb.clk_d14 ;
 wire \u_skew_usb.clk_d15 ;
 wire \u_skew_usb.clk_d2 ;
 wire \u_skew_usb.clk_d3 ;
 wire \u_skew_usb.clk_d4 ;
 wire \u_skew_usb.clk_d5 ;
 wire \u_skew_usb.clk_d6 ;
 wire \u_skew_usb.clk_d7 ;
 wire \u_skew_usb.clk_d8 ;
 wire \u_skew_usb.clk_d9 ;
 wire \u_skew_usb.clk_inbuf ;
 wire \u_skew_usb.clkbuf_1.X1 ;
 wire \u_skew_usb.clkbuf_1.X2 ;
 wire \u_skew_usb.clkbuf_1.X3 ;
 wire \u_skew_usb.clkbuf_10.X1 ;
 wire \u_skew_usb.clkbuf_10.X2 ;
 wire \u_skew_usb.clkbuf_10.X3 ;
 wire \u_skew_usb.clkbuf_11.X1 ;
 wire \u_skew_usb.clkbuf_11.X2 ;
 wire \u_skew_usb.clkbuf_11.X3 ;
 wire \u_skew_usb.clkbuf_12.X1 ;
 wire \u_skew_usb.clkbuf_12.X2 ;
 wire \u_skew_usb.clkbuf_12.X3 ;
 wire \u_skew_usb.clkbuf_13.X1 ;
 wire \u_skew_usb.clkbuf_13.X2 ;
 wire \u_skew_usb.clkbuf_13.X3 ;
 wire \u_skew_usb.clkbuf_14.X1 ;
 wire \u_skew_usb.clkbuf_14.X2 ;
 wire \u_skew_usb.clkbuf_14.X3 ;
 wire \u_skew_usb.clkbuf_15.X1 ;
 wire \u_skew_usb.clkbuf_15.X2 ;
 wire \u_skew_usb.clkbuf_15.X3 ;
 wire \u_skew_usb.clkbuf_2.X1 ;
 wire \u_skew_usb.clkbuf_2.X2 ;
 wire \u_skew_usb.clkbuf_2.X3 ;
 wire \u_skew_usb.clkbuf_3.X1 ;
 wire \u_skew_usb.clkbuf_3.X2 ;
 wire \u_skew_usb.clkbuf_3.X3 ;
 wire \u_skew_usb.clkbuf_4.X1 ;
 wire \u_skew_usb.clkbuf_4.X2 ;
 wire \u_skew_usb.clkbuf_4.X3 ;
 wire \u_skew_usb.clkbuf_5.X1 ;
 wire \u_skew_usb.clkbuf_5.X2 ;
 wire \u_skew_usb.clkbuf_5.X3 ;
 wire \u_skew_usb.clkbuf_6.X1 ;
 wire \u_skew_usb.clkbuf_6.X2 ;
 wire \u_skew_usb.clkbuf_6.X3 ;
 wire \u_skew_usb.clkbuf_7.X1 ;
 wire \u_skew_usb.clkbuf_7.X2 ;
 wire \u_skew_usb.clkbuf_7.X3 ;
 wire \u_skew_usb.clkbuf_8.X1 ;
 wire \u_skew_usb.clkbuf_8.X2 ;
 wire \u_skew_usb.clkbuf_8.X3 ;
 wire \u_skew_usb.clkbuf_9.X1 ;
 wire \u_skew_usb.clkbuf_9.X2 ;
 wire \u_skew_usb.clkbuf_9.X3 ;
 wire \u_skew_usb.d00 ;
 wire \u_skew_usb.d01 ;
 wire \u_skew_usb.d02 ;
 wire \u_skew_usb.d03 ;
 wire \u_skew_usb.d04 ;
 wire \u_skew_usb.d05 ;
 wire \u_skew_usb.d06 ;
 wire \u_skew_usb.d07 ;
 wire \u_skew_usb.d10 ;
 wire \u_skew_usb.d11 ;
 wire \u_skew_usb.d12 ;
 wire \u_skew_usb.d13 ;
 wire \u_skew_usb.d20 ;
 wire \u_skew_usb.d21 ;
 wire \u_skew_usb.d30 ;
 wire \u_skew_usb.in0 ;
 wire \u_skew_usb.in1 ;
 wire \u_skew_usb.in10 ;
 wire \u_skew_usb.in11 ;
 wire \u_skew_usb.in12 ;
 wire \u_skew_usb.in13 ;
 wire \u_skew_usb.in14 ;
 wire \u_skew_usb.in15 ;
 wire \u_skew_usb.in2 ;
 wire \u_skew_usb.in3 ;
 wire \u_skew_usb.in4 ;
 wire \u_skew_usb.in5 ;
 wire \u_skew_usb.in6 ;
 wire \u_skew_usb.in7 ;
 wire \u_skew_usb.in8 ;
 wire \u_skew_usb.in9 ;
 wire \u_usb_host.reg_ack ;
 wire \u_usb_host.reg_addr[0] ;
 wire \u_usb_host.reg_addr[1] ;
 wire \u_usb_host.reg_addr[2] ;
 wire \u_usb_host.reg_addr[3] ;
 wire \u_usb_host.reg_addr[4] ;
 wire \u_usb_host.reg_addr[5] ;
 wire \u_usb_host.reg_cs ;
 wire \u_usb_host.reg_rdata[0] ;
 wire \u_usb_host.reg_rdata[10] ;
 wire \u_usb_host.reg_rdata[11] ;
 wire \u_usb_host.reg_rdata[12] ;
 wire \u_usb_host.reg_rdata[13] ;
 wire \u_usb_host.reg_rdata[14] ;
 wire \u_usb_host.reg_rdata[15] ;
 wire \u_usb_host.reg_rdata[16] ;
 wire \u_usb_host.reg_rdata[17] ;
 wire \u_usb_host.reg_rdata[18] ;
 wire \u_usb_host.reg_rdata[19] ;
 wire \u_usb_host.reg_rdata[1] ;
 wire \u_usb_host.reg_rdata[20] ;
 wire \u_usb_host.reg_rdata[21] ;
 wire \u_usb_host.reg_rdata[22] ;
 wire \u_usb_host.reg_rdata[23] ;
 wire \u_usb_host.reg_rdata[24] ;
 wire \u_usb_host.reg_rdata[25] ;
 wire \u_usb_host.reg_rdata[26] ;
 wire \u_usb_host.reg_rdata[27] ;
 wire \u_usb_host.reg_rdata[28] ;
 wire \u_usb_host.reg_rdata[29] ;
 wire \u_usb_host.reg_rdata[2] ;
 wire \u_usb_host.reg_rdata[30] ;
 wire \u_usb_host.reg_rdata[31] ;
 wire \u_usb_host.reg_rdata[3] ;
 wire \u_usb_host.reg_rdata[4] ;
 wire \u_usb_host.reg_rdata[5] ;
 wire \u_usb_host.reg_rdata[6] ;
 wire \u_usb_host.reg_rdata[7] ;
 wire \u_usb_host.reg_rdata[8] ;
 wire \u_usb_host.reg_rdata[9] ;
 wire \u_usb_host.reg_wdata[0] ;
 wire \u_usb_host.reg_wdata[10] ;
 wire \u_usb_host.reg_wdata[11] ;
 wire \u_usb_host.reg_wdata[12] ;
 wire \u_usb_host.reg_wdata[13] ;
 wire \u_usb_host.reg_wdata[14] ;
 wire \u_usb_host.reg_wdata[15] ;
 wire \u_usb_host.reg_wdata[16] ;
 wire \u_usb_host.reg_wdata[17] ;
 wire \u_usb_host.reg_wdata[18] ;
 wire \u_usb_host.reg_wdata[19] ;
 wire \u_usb_host.reg_wdata[1] ;
 wire \u_usb_host.reg_wdata[20] ;
 wire \u_usb_host.reg_wdata[21] ;
 wire \u_usb_host.reg_wdata[22] ;
 wire \u_usb_host.reg_wdata[23] ;
 wire \u_usb_host.reg_wdata[28] ;
 wire \u_usb_host.reg_wdata[29] ;
 wire \u_usb_host.reg_wdata[2] ;
 wire \u_usb_host.reg_wdata[30] ;
 wire \u_usb_host.reg_wdata[31] ;
 wire \u_usb_host.reg_wdata[3] ;
 wire \u_usb_host.reg_wdata[4] ;
 wire \u_usb_host.reg_wdata[5] ;
 wire \u_usb_host.reg_wdata[6] ;
 wire \u_usb_host.reg_wdata[7] ;
 wire \u_usb_host.reg_wdata[8] ;
 wire \u_usb_host.reg_wdata[9] ;
 wire \u_usb_host.reg_wr ;
 wire \u_usb_host.u_async_wb.PendingRd ;
 wire \u_usb_host.u_async_wb._00_ ;
 wire \u_usb_host.u_async_wb._01_ ;
 wire \u_usb_host.u_async_wb._02_ ;
 wire \u_usb_host.u_async_wb._03_ ;
 wire \u_usb_host.u_async_wb._04_ ;
 wire \u_usb_host.u_async_wb._05_ ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_afull ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_en ;
 wire \u_usb_host.u_async_wb.m_cmd_wr_full ;
 wire \u_usb_host.u_async_wb.m_resp_rd_empty ;
 wire \u_usb_host.u_async_wb.m_resp_rd_en ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[10] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[11] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[12] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[13] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[14] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[15] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[16] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[17] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[18] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[19] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[20] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[21] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[22] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[23] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[24] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[25] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[26] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[27] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[32] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[33] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[34] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[35] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[36] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[37] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[38] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[39] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[40] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[41] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[42] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[4] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[5] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[6] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[7] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[8] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_data[9] ;
 wire \u_usb_host.u_async_wb.s_cmd_rd_empty ;
 wire \u_usb_host.u_async_wb.s_resp_wr_en ;
 wire \u_usb_host.u_async_wb.s_resp_wr_full ;
 wire \u_usb_host.u_async_wb.u_cmd_if._000_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._001_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._002_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._003_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._004_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._005_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._006_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._007_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._008_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._009_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._010_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._011_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._012_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._013_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._014_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._015_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._016_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._017_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._018_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._019_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._020_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._021_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._022_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._023_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._024_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._025_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._026_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._027_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._030_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._031_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._033_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._034_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._035_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._036_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._037_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._038_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._039_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._040_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._041_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if._042_ ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ;
 wire \u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ;
 wire \u_usb_host.u_async_wb.u_resp_if._000_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._001_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._002_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._003_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._004_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._005_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._006_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._007_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._008_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._009_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._010_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._011_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._012_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._013_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._014_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._015_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._016_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._017_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._018_ ;
 wire \u_usb_host.u_async_wb.u_resp_if._019_ ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[0][9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.mem[1][9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[10] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[11] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[12] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[13] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[14] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[15] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[16] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[17] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[18] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[19] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[20] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[21] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[22] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[23] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[24] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[25] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[26] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[27] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[28] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[29] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[2] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[30] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[31] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[3] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[4] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[5] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[6] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[7] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[8] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_data[9] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ;
 wire \u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ;
 wire \u_usb_host.u_async_wb.wbm_cyc_i ;
 wire \u_usb_host.u_async_wb.wbs_ack_f ;
 wire \u_usb_host.u_async_wb.wbs_cyc_o ;
 wire \u_usb_host.u_core._000_ ;
 wire \u_usb_host.u_core._001_ ;
 wire \u_usb_host.u_core._002_ ;
 wire \u_usb_host.u_core._003_ ;
 wire \u_usb_host.u_core._004_ ;
 wire \u_usb_host.u_core._005_ ;
 wire \u_usb_host.u_core._006_ ;
 wire \u_usb_host.u_core._007_ ;
 wire \u_usb_host.u_core._008_ ;
 wire \u_usb_host.u_core._009_ ;
 wire \u_usb_host.u_core._010_ ;
 wire \u_usb_host.u_core._011_ ;
 wire \u_usb_host.u_core._012_ ;
 wire \u_usb_host.u_core._013_ ;
 wire \u_usb_host.u_core._014_ ;
 wire \u_usb_host.u_core._015_ ;
 wire \u_usb_host.u_core._016_ ;
 wire \u_usb_host.u_core._017_ ;
 wire \u_usb_host.u_core._018_ ;
 wire \u_usb_host.u_core._019_ ;
 wire \u_usb_host.u_core._020_ ;
 wire \u_usb_host.u_core._021_ ;
 wire \u_usb_host.u_core._022_ ;
 wire \u_usb_host.u_core._023_ ;
 wire \u_usb_host.u_core._024_ ;
 wire \u_usb_host.u_core._025_ ;
 wire \u_usb_host.u_core._026_ ;
 wire \u_usb_host.u_core._027_ ;
 wire \u_usb_host.u_core._028_ ;
 wire \u_usb_host.u_core._029_ ;
 wire \u_usb_host.u_core._030_ ;
 wire \u_usb_host.u_core._031_ ;
 wire \u_usb_host.u_core._032_ ;
 wire \u_usb_host.u_core._033_ ;
 wire \u_usb_host.u_core._034_ ;
 wire \u_usb_host.u_core._035_ ;
 wire \u_usb_host.u_core._036_ ;
 wire \u_usb_host.u_core._037_ ;
 wire \u_usb_host.u_core._038_ ;
 wire \u_usb_host.u_core._039_ ;
 wire \u_usb_host.u_core._040_ ;
 wire \u_usb_host.u_core._041_ ;
 wire \u_usb_host.u_core._042_ ;
 wire \u_usb_host.u_core._043_ ;
 wire \u_usb_host.u_core._044_ ;
 wire \u_usb_host.u_core._045_ ;
 wire \u_usb_host.u_core._046_ ;
 wire \u_usb_host.u_core._047_ ;
 wire \u_usb_host.u_core._048_ ;
 wire \u_usb_host.u_core._049_ ;
 wire \u_usb_host.u_core._050_ ;
 wire \u_usb_host.u_core._051_ ;
 wire \u_usb_host.u_core._052_ ;
 wire \u_usb_host.u_core._053_ ;
 wire \u_usb_host.u_core._054_ ;
 wire \u_usb_host.u_core._055_ ;
 wire \u_usb_host.u_core._056_ ;
 wire \u_usb_host.u_core._057_ ;
 wire \u_usb_host.u_core._058_ ;
 wire \u_usb_host.u_core._059_ ;
 wire \u_usb_host.u_core._060_ ;
 wire \u_usb_host.u_core._061_ ;
 wire \u_usb_host.u_core._062_ ;
 wire \u_usb_host.u_core._063_ ;
 wire \u_usb_host.u_core._064_ ;
 wire \u_usb_host.u_core._065_ ;
 wire \u_usb_host.u_core._066_ ;
 wire \u_usb_host.u_core._067_ ;
 wire \u_usb_host.u_core._068_ ;
 wire \u_usb_host.u_core._069_ ;
 wire \u_usb_host.u_core._070_ ;
 wire \u_usb_host.u_core._071_ ;
 wire \u_usb_host.u_core._072_ ;
 wire \u_usb_host.u_core._073_ ;
 wire \u_usb_host.u_core._074_ ;
 wire \u_usb_host.u_core._075_ ;
 wire \u_usb_host.u_core._076_ ;
 wire \u_usb_host.u_core._077_ ;
 wire \u_usb_host.u_core._078_ ;
 wire \u_usb_host.u_core._079_ ;
 wire \u_usb_host.u_core._080_ ;
 wire \u_usb_host.u_core._081_ ;
 wire \u_usb_host.u_core._082_ ;
 wire \u_usb_host.u_core._083_ ;
 wire \u_usb_host.u_core._084_ ;
 wire \u_usb_host.u_core._085_ ;
 wire \u_usb_host.u_core._086_ ;
 wire \u_usb_host.u_core._087_ ;
 wire \u_usb_host.u_core._088_ ;
 wire \u_usb_host.u_core._089_ ;
 wire \u_usb_host.u_core._090_ ;
 wire \u_usb_host.u_core._091_ ;
 wire \u_usb_host.u_core._092_ ;
 wire \u_usb_host.u_core._093_ ;
 wire \u_usb_host.u_core._094_ ;
 wire \u_usb_host.u_core._095_ ;
 wire \u_usb_host.u_core._096_ ;
 wire \u_usb_host.u_core._097_ ;
 wire \u_usb_host.u_core._098_ ;
 wire \u_usb_host.u_core._099_ ;
 wire \u_usb_host.u_core._100_ ;
 wire \u_usb_host.u_core._101_ ;
 wire \u_usb_host.u_core._102_ ;
 wire \u_usb_host.u_core._103_ ;
 wire \u_usb_host.u_core._104_ ;
 wire \u_usb_host.u_core._105_ ;
 wire \u_usb_host.u_core._106_ ;
 wire \u_usb_host.u_core._107_ ;
 wire \u_usb_host.u_core._108_ ;
 wire \u_usb_host.u_core._109_ ;
 wire \u_usb_host.u_core._110_ ;
 wire \u_usb_host.u_core._111_ ;
 wire \u_usb_host.u_core._112_ ;
 wire \u_usb_host.u_core._113_ ;
 wire \u_usb_host.u_core._114_ ;
 wire \u_usb_host.u_core._115_ ;
 wire \u_usb_host.u_core._116_ ;
 wire \u_usb_host.u_core._117_ ;
 wire \u_usb_host.u_core._118_ ;
 wire \u_usb_host.u_core._119_ ;
 wire \u_usb_host.u_core._120_ ;
 wire \u_usb_host.u_core._121_ ;
 wire \u_usb_host.u_core._122_ ;
 wire \u_usb_host.u_core._123_ ;
 wire \u_usb_host.u_core._124_ ;
 wire \u_usb_host.u_core._125_ ;
 wire \u_usb_host.u_core._126_ ;
 wire \u_usb_host.u_core._127_ ;
 wire \u_usb_host.u_core._128_ ;
 wire \u_usb_host.u_core._129_ ;
 wire \u_usb_host.u_core._130_ ;
 wire \u_usb_host.u_core._131_ ;
 wire \u_usb_host.u_core._132_ ;
 wire \u_usb_host.u_core._133_ ;
 wire \u_usb_host.u_core._134_ ;
 wire \u_usb_host.u_core._135_ ;
 wire \u_usb_host.u_core._136_ ;
 wire \u_usb_host.u_core._137_ ;
 wire \u_usb_host.u_core._138_ ;
 wire \u_usb_host.u_core._139_ ;
 wire \u_usb_host.u_core._140_ ;
 wire \u_usb_host.u_core._141_ ;
 wire \u_usb_host.u_core._142_ ;
 wire \u_usb_host.u_core._143_ ;
 wire \u_usb_host.u_core._144_ ;
 wire \u_usb_host.u_core._145_ ;
 wire \u_usb_host.u_core._146_ ;
 wire \u_usb_host.u_core._147_ ;
 wire \u_usb_host.u_core._148_ ;
 wire \u_usb_host.u_core._149_ ;
 wire \u_usb_host.u_core._150_ ;
 wire \u_usb_host.u_core._151_ ;
 wire \u_usb_host.u_core._152_ ;
 wire \u_usb_host.u_core._153_ ;
 wire \u_usb_host.u_core._154_ ;
 wire \u_usb_host.u_core._155_ ;
 wire \u_usb_host.u_core._156_ ;
 wire \u_usb_host.u_core._157_ ;
 wire \u_usb_host.u_core._158_ ;
 wire \u_usb_host.u_core._159_ ;
 wire \u_usb_host.u_core._160_ ;
 wire \u_usb_host.u_core._161_ ;
 wire \u_usb_host.u_core._162_ ;
 wire \u_usb_host.u_core._163_ ;
 wire \u_usb_host.u_core._164_ ;
 wire \u_usb_host.u_core._165_ ;
 wire \u_usb_host.u_core._166_ ;
 wire \u_usb_host.u_core._167_ ;
 wire \u_usb_host.u_core._168_ ;
 wire \u_usb_host.u_core._169_ ;
 wire \u_usb_host.u_core._170_ ;
 wire \u_usb_host.u_core._171_ ;
 wire \u_usb_host.u_core._172_ ;
 wire \u_usb_host.u_core._173_ ;
 wire \u_usb_host.u_core._174_ ;
 wire \u_usb_host.u_core._175_ ;
 wire \u_usb_host.u_core._176_ ;
 wire \u_usb_host.u_core._177_ ;
 wire \u_usb_host.u_core._178_ ;
 wire \u_usb_host.u_core._179_ ;
 wire \u_usb_host.u_core._180_ ;
 wire \u_usb_host.u_core._181_ ;
 wire \u_usb_host.u_core._182_ ;
 wire \u_usb_host.u_core._183_ ;
 wire \u_usb_host.u_core._184_ ;
 wire \u_usb_host.u_core._185_ ;
 wire \u_usb_host.u_core._186_ ;
 wire \u_usb_host.u_core._187_ ;
 wire \u_usb_host.u_core._188_ ;
 wire \u_usb_host.u_core._189_ ;
 wire \u_usb_host.u_core._190_ ;
 wire \u_usb_host.u_core._191_ ;
 wire \u_usb_host.u_core._192_ ;
 wire \u_usb_host.u_core._193_ ;
 wire \u_usb_host.u_core._194_ ;
 wire \u_usb_host.u_core._195_ ;
 wire \u_usb_host.u_core._196_ ;
 wire \u_usb_host.u_core._197_ ;
 wire \u_usb_host.u_core._198_ ;
 wire \u_usb_host.u_core._199_ ;
 wire \u_usb_host.u_core._200_ ;
 wire \u_usb_host.u_core._201_ ;
 wire \u_usb_host.u_core._202_ ;
 wire \u_usb_host.u_core.cfg_wr ;
 wire \u_usb_host.u_core.device_det_q ;
 wire \u_usb_host.u_core.err_cond_q ;
 wire \u_usb_host.u_core.fifo_flush_q ;
 wire \u_usb_host.u_core.fifo_rx_data_w[0] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[1] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[2] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[3] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[4] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[5] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[6] ;
 wire \u_usb_host.u_core.fifo_rx_data_w[7] ;
 wire \u_usb_host.u_core.fifo_rx_push_w ;
 wire \u_usb_host.u_core.fifo_tx_data_w[0] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[1] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[2] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[3] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[4] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[5] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[6] ;
 wire \u_usb_host.u_core.fifo_tx_data_w[7] ;
 wire \u_usb_host.u_core.fifo_tx_pop_w ;
 wire \u_usb_host.u_core.in_transfer_q ;
 wire \u_usb_host.u_core.intr_done_q ;
 wire \u_usb_host.u_core.intr_err_q ;
 wire \u_usb_host.u_core.intr_sof_q ;
 wire \u_usb_host.u_core.reg_rdata_r[0] ;
 wire \u_usb_host.u_core.reg_rdata_r[10] ;
 wire \u_usb_host.u_core.reg_rdata_r[11] ;
 wire \u_usb_host.u_core.reg_rdata_r[12] ;
 wire \u_usb_host.u_core.reg_rdata_r[13] ;
 wire \u_usb_host.u_core.reg_rdata_r[14] ;
 wire \u_usb_host.u_core.reg_rdata_r[15] ;
 wire \u_usb_host.u_core.reg_rdata_r[16] ;
 wire \u_usb_host.u_core.reg_rdata_r[17] ;
 wire \u_usb_host.u_core.reg_rdata_r[18] ;
 wire \u_usb_host.u_core.reg_rdata_r[19] ;
 wire \u_usb_host.u_core.reg_rdata_r[1] ;
 wire \u_usb_host.u_core.reg_rdata_r[20] ;
 wire \u_usb_host.u_core.reg_rdata_r[21] ;
 wire \u_usb_host.u_core.reg_rdata_r[22] ;
 wire \u_usb_host.u_core.reg_rdata_r[23] ;
 wire \u_usb_host.u_core.reg_rdata_r[24] ;
 wire \u_usb_host.u_core.reg_rdata_r[25] ;
 wire \u_usb_host.u_core.reg_rdata_r[26] ;
 wire \u_usb_host.u_core.reg_rdata_r[27] ;
 wire \u_usb_host.u_core.reg_rdata_r[28] ;
 wire \u_usb_host.u_core.reg_rdata_r[29] ;
 wire \u_usb_host.u_core.reg_rdata_r[2] ;
 wire \u_usb_host.u_core.reg_rdata_r[30] ;
 wire \u_usb_host.u_core.reg_rdata_r[31] ;
 wire \u_usb_host.u_core.reg_rdata_r[3] ;
 wire \u_usb_host.u_core.reg_rdata_r[4] ;
 wire \u_usb_host.u_core.reg_rdata_r[5] ;
 wire \u_usb_host.u_core.reg_rdata_r[6] ;
 wire \u_usb_host.u_core.reg_rdata_r[7] ;
 wire \u_usb_host.u_core.reg_rdata_r[8] ;
 wire \u_usb_host.u_core.reg_rdata_r[9] ;
 wire \u_usb_host.u_core.resp_expected_q ;
 wire \u_usb_host.u_core.send_sof_w ;
 wire \u_usb_host.u_core.sof_irq_q ;
 wire \u_usb_host.u_core.sof_time_q[0] ;
 wire \u_usb_host.u_core.sof_time_q[10] ;
 wire \u_usb_host.u_core.sof_time_q[11] ;
 wire \u_usb_host.u_core.sof_time_q[12] ;
 wire \u_usb_host.u_core.sof_time_q[13] ;
 wire \u_usb_host.u_core.sof_time_q[14] ;
 wire \u_usb_host.u_core.sof_time_q[15] ;
 wire \u_usb_host.u_core.sof_time_q[1] ;
 wire \u_usb_host.u_core.sof_time_q[2] ;
 wire \u_usb_host.u_core.sof_time_q[3] ;
 wire \u_usb_host.u_core.sof_time_q[4] ;
 wire \u_usb_host.u_core.sof_time_q[5] ;
 wire \u_usb_host.u_core.sof_time_q[6] ;
 wire \u_usb_host.u_core.sof_time_q[7] ;
 wire \u_usb_host.u_core.sof_time_q[8] ;
 wire \u_usb_host.u_core.sof_time_q[9] ;
 wire \u_usb_host.u_core.sof_transfer_q ;
 wire \u_usb_host.u_core.sof_value_q[0] ;
 wire \u_usb_host.u_core.sof_value_q[10] ;
 wire \u_usb_host.u_core.sof_value_q[1] ;
 wire \u_usb_host.u_core.sof_value_q[2] ;
 wire \u_usb_host.u_core.sof_value_q[3] ;
 wire \u_usb_host.u_core.sof_value_q[4] ;
 wire \u_usb_host.u_core.sof_value_q[5] ;
 wire \u_usb_host.u_core.sof_value_q[6] ;
 wire \u_usb_host.u_core.sof_value_q[7] ;
 wire \u_usb_host.u_core.sof_value_q[8] ;
 wire \u_usb_host.u_core.sof_value_q[9] ;
 wire \u_usb_host.u_core.status_crc_err_w ;
 wire \u_usb_host.u_core.status_response_w[0] ;
 wire \u_usb_host.u_core.status_response_w[1] ;
 wire \u_usb_host.u_core.status_response_w[2] ;
 wire \u_usb_host.u_core.status_response_w[3] ;
 wire \u_usb_host.u_core.status_response_w[4] ;
 wire \u_usb_host.u_core.status_response_w[5] ;
 wire \u_usb_host.u_core.status_response_w[6] ;
 wire \u_usb_host.u_core.status_response_w[7] ;
 wire \u_usb_host.u_core.status_rx_count_w[0] ;
 wire \u_usb_host.u_core.status_rx_count_w[10] ;
 wire \u_usb_host.u_core.status_rx_count_w[11] ;
 wire \u_usb_host.u_core.status_rx_count_w[12] ;
 wire \u_usb_host.u_core.status_rx_count_w[13] ;
 wire \u_usb_host.u_core.status_rx_count_w[14] ;
 wire \u_usb_host.u_core.status_rx_count_w[15] ;
 wire \u_usb_host.u_core.status_rx_count_w[1] ;
 wire \u_usb_host.u_core.status_rx_count_w[2] ;
 wire \u_usb_host.u_core.status_rx_count_w[3] ;
 wire \u_usb_host.u_core.status_rx_count_w[4] ;
 wire \u_usb_host.u_core.status_rx_count_w[5] ;
 wire \u_usb_host.u_core.status_rx_count_w[6] ;
 wire \u_usb_host.u_core.status_rx_count_w[7] ;
 wire \u_usb_host.u_core.status_rx_count_w[8] ;
 wire \u_usb_host.u_core.status_rx_count_w[9] ;
 wire \u_usb_host.u_core.status_rx_done_w ;
 wire \u_usb_host.u_core.status_sie_idle_w ;
 wire \u_usb_host.u_core.status_timeout_w ;
 wire \u_usb_host.u_core.status_tx_done_w ;
 wire \u_usb_host.u_core.token_dev_w[0] ;
 wire \u_usb_host.u_core.token_dev_w[1] ;
 wire \u_usb_host.u_core.token_dev_w[2] ;
 wire \u_usb_host.u_core.token_dev_w[3] ;
 wire \u_usb_host.u_core.token_dev_w[4] ;
 wire \u_usb_host.u_core.token_dev_w[5] ;
 wire \u_usb_host.u_core.token_dev_w[6] ;
 wire \u_usb_host.u_core.token_ep_w[0] ;
 wire \u_usb_host.u_core.token_ep_w[1] ;
 wire \u_usb_host.u_core.token_ep_w[2] ;
 wire \u_usb_host.u_core.token_ep_w[3] ;
 wire \u_usb_host.u_core.token_pid_w[0] ;
 wire \u_usb_host.u_core.token_pid_w[1] ;
 wire \u_usb_host.u_core.token_pid_w[2] ;
 wire \u_usb_host.u_core.token_pid_w[3] ;
 wire \u_usb_host.u_core.token_pid_w[4] ;
 wire \u_usb_host.u_core.token_pid_w[5] ;
 wire \u_usb_host.u_core.token_pid_w[6] ;
 wire \u_usb_host.u_core.token_pid_w[7] ;
 wire \u_usb_host.u_core.transfer_ack_w ;
 wire \u_usb_host.u_core.transfer_start_q ;
 wire \u_usb_host.u_core.u_fifo_rx._0000_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0001_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0002_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0003_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0004_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0005_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0006_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0007_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0008_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0009_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0010_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0011_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0012_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0013_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0014_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0015_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0016_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0017_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0018_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0019_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0020_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0021_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0022_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0023_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0024_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0025_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0026_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0027_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0028_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0029_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0030_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0031_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0032_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0033_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0034_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0035_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0036_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0037_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0038_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0039_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0040_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0041_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0042_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0043_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0044_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0045_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0046_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0047_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0048_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0049_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0050_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0051_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0052_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0053_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0054_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0055_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0056_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0057_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0058_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0059_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0060_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0061_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0062_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0063_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0064_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0065_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0066_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0067_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0068_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0069_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0070_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0071_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0072_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0073_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0074_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0075_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0076_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0077_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0078_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0079_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0080_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0081_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0082_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0083_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0084_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0085_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0086_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0087_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0088_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0089_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0090_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0091_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0092_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0093_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0094_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0095_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0096_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0097_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0098_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0099_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0100_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0101_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0102_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0103_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0104_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0105_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0106_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0107_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0108_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0109_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0110_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0111_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0112_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0113_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0114_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0115_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0116_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0117_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0118_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0119_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0120_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0121_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0122_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0123_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0124_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0125_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0126_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0127_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0128_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0129_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0130_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0131_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0132_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0133_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0134_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0135_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0136_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0137_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0138_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0139_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0140_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0141_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0142_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0143_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0144_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0145_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0146_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0147_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0148_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0149_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0150_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0151_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0152_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0153_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0154_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0155_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0156_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0157_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0158_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0159_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0160_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0161_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0162_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0163_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0164_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0165_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0166_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0167_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0168_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0169_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0170_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0171_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0172_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0173_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0174_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0175_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0176_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0177_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0178_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0179_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0180_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0181_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0182_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0183_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0184_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0185_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0186_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0187_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0188_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0189_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0190_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0191_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0192_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0193_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0194_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0195_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0196_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0197_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0198_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0199_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0200_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0201_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0202_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0203_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0204_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0205_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0206_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0207_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0208_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0209_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0210_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0211_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0212_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0213_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0214_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0215_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0216_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0217_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0218_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0219_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0220_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0221_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0222_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0223_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0224_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0225_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0226_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0227_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0228_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0229_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0230_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0231_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0232_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0233_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0234_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0235_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0236_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0237_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0238_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0239_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0240_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0241_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0242_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0243_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0244_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0245_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0246_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0247_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0248_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0249_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0250_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0251_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0252_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0253_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0254_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0255_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0256_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0257_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0258_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0259_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0260_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0261_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0262_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0263_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0264_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0265_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0266_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0267_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0268_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0269_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0270_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0271_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0272_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0273_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0274_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0275_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0276_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0277_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0278_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0279_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0280_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0281_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0282_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0283_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0284_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0285_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0286_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0287_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0288_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0289_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0290_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0291_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0292_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0293_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0294_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0295_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0296_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0297_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0298_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0299_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0300_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0301_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0302_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0303_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0304_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0305_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0306_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0307_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0308_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0309_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0310_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0311_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0312_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0313_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0314_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0315_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0316_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0317_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0318_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0319_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0320_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0321_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0322_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0323_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0324_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0325_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0326_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0327_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0328_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0329_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0330_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0331_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0332_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0333_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0334_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0335_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0336_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0337_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0338_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0339_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0340_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0341_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0342_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0343_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0344_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0345_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0346_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0347_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0348_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0349_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0350_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0351_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0352_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0353_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0354_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0355_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0356_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0357_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0358_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0359_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0360_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0361_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0362_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0363_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0364_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0365_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0366_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0367_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0368_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0369_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0370_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0371_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0372_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0373_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0374_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0375_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0376_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0377_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0378_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0379_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0380_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0381_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0382_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0383_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0384_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0385_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0386_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0387_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0388_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0389_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0390_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0391_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0392_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0393_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0394_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0395_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0396_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0397_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0398_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0399_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0400_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0401_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0402_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0403_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0404_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0405_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0406_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0407_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0408_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0409_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0410_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0411_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0412_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0413_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0414_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0415_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0416_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0417_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0418_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0419_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0420_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0421_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0422_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0423_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0424_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0425_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0426_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0427_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0428_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0429_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0430_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0431_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0432_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0433_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0434_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0435_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0436_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0437_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0438_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0439_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0440_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0441_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0442_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0443_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0444_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0445_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0446_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0447_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0448_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0449_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0450_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0451_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0452_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0453_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0454_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0455_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0456_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0457_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0458_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0459_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0460_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0461_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0462_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0463_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0464_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0465_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0466_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0467_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0468_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0469_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0470_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0471_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0472_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0473_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0474_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0475_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0476_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0477_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0478_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0479_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0480_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0481_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0482_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0483_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0484_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0485_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0486_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0487_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0488_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0489_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0490_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0491_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0492_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0493_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0494_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0495_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0496_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0497_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0498_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0499_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0500_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0501_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0502_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0503_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0504_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0505_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0506_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0507_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0508_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0509_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0510_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0511_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0512_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0513_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0514_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0515_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0516_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0517_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0518_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0519_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0520_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0521_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0522_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0523_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0524_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0525_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0526_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0527_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0528_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0529_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0530_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0531_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0532_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0533_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0534_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0535_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0536_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0537_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0538_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0539_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0540_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0541_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0542_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0543_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0544_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0545_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0546_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0547_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0548_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0549_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0550_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0551_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0552_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0553_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0554_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0555_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0556_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0557_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0558_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0559_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0560_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0561_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0562_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0563_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0564_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0565_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0566_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0567_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0568_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0569_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0570_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0571_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0572_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0573_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0574_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0575_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0576_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0577_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0578_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0579_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0580_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0581_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0582_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0583_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0584_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0585_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0586_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0587_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0588_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0589_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0590_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0591_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0592_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0593_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0594_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0595_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0596_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0597_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0598_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0599_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0600_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0601_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0602_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0603_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0604_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0605_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0606_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0607_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0608_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0609_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0610_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0611_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0612_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0613_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0614_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0615_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0616_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0617_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0618_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0619_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0620_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0621_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0622_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0623_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0624_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0625_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0626_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0627_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0628_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0629_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0630_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0631_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0632_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0633_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0634_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0635_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0636_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0637_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0638_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0639_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0640_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0641_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0642_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0643_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0644_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0645_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0646_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0647_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0648_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0649_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0650_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0651_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0652_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0653_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0654_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0655_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0656_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0657_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0658_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0659_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0660_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0661_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0662_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0663_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0664_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0665_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0666_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0667_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0668_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0669_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0670_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0671_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0672_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0673_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0674_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0675_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0676_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0677_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0678_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0679_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0680_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0681_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0682_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0683_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0684_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0685_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0686_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0687_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0688_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0689_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0690_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0691_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0692_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0693_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0694_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0695_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0696_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0697_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0698_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0699_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0700_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0701_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0702_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0703_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0704_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0705_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0706_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0707_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0708_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0709_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0710_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0711_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0712_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0713_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0714_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0715_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0716_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0717_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0718_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0719_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0720_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0721_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0722_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0723_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0724_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0725_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0726_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0727_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0728_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0729_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0730_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0731_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0732_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0733_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0734_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0735_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0736_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0737_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0738_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0739_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0740_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0741_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0742_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0743_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0744_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0745_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0746_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0747_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0748_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0749_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0750_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0751_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0752_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0753_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0754_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0755_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0756_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0757_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0758_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0759_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0760_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0761_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0762_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0763_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0764_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0765_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0766_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0767_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0768_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0769_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0770_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0771_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0772_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0773_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0774_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0775_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0776_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0777_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0778_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0779_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0780_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0781_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0782_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0783_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0784_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0785_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0786_ ;
 wire \u_usb_host.u_core.u_fifo_rx._0787_ ;
 wire \u_usb_host.u_core.u_fifo_rx.count[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.count[6] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[6] ;
 wire \u_usb_host.u_core.u_fifo_rx.data_o[7] ;
 wire \u_usb_host.u_core.u_fifo_rx.pop_i ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[0][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[10][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[11][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[12][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[13][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[14][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[15][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[16][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[17][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[18][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[19][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[1][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[20][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[21][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[22][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[23][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[24][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[25][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[26][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[27][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[28][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[29][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[2][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[30][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[31][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[32][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[33][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[34][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[35][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[36][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[37][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[38][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[39][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[3][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[40][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[41][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[42][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[43][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[44][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[45][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[46][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[47][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[48][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[49][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[4][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[50][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[51][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[52][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[53][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[54][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[55][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[56][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[57][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[58][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[59][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[5][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[60][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[61][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[62][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[63][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[6][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[7][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[8][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][0] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][1] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][2] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][3] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][4] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][5] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][6] ;
 wire \u_usb_host.u_core.u_fifo_rx.ram[9][7] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ;
 wire \u_usb_host.u_core.u_fifo_tx._0000_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0001_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0002_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0003_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0004_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0005_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0006_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0007_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0008_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0009_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0010_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0011_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0012_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0013_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0014_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0015_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0016_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0017_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0018_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0019_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0020_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0021_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0022_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0023_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0024_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0025_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0026_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0027_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0028_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0029_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0030_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0031_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0032_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0033_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0034_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0035_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0036_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0037_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0038_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0039_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0040_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0041_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0042_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0043_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0044_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0045_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0046_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0047_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0048_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0049_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0050_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0051_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0052_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0053_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0054_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0055_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0056_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0057_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0058_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0059_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0060_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0061_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0062_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0063_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0064_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0065_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0066_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0067_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0068_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0069_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0070_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0071_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0072_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0073_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0074_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0075_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0076_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0077_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0078_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0079_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0080_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0081_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0082_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0083_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0084_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0085_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0086_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0087_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0088_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0089_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0090_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0091_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0092_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0093_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0094_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0095_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0096_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0097_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0098_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0099_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0100_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0101_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0102_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0103_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0104_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0105_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0106_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0107_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0108_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0109_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0110_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0111_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0112_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0113_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0114_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0115_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0116_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0117_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0118_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0119_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0120_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0121_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0122_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0123_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0124_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0125_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0126_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0127_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0128_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0129_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0130_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0131_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0132_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0133_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0134_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0135_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0136_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0137_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0138_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0139_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0140_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0141_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0142_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0143_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0144_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0145_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0146_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0147_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0148_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0149_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0150_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0151_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0152_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0153_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0154_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0155_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0156_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0157_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0158_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0159_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0160_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0161_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0162_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0163_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0164_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0165_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0166_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0167_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0168_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0169_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0170_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0171_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0172_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0173_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0174_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0175_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0176_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0177_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0178_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0179_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0180_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0181_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0182_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0183_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0184_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0185_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0186_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0187_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0188_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0189_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0190_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0191_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0192_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0193_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0194_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0195_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0196_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0197_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0198_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0199_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0200_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0201_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0202_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0203_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0204_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0205_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0206_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0207_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0208_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0209_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0210_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0211_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0212_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0213_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0214_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0215_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0216_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0217_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0218_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0219_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0220_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0221_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0222_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0223_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0224_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0225_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0226_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0227_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0228_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0229_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0230_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0231_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0232_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0233_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0234_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0235_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0236_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0237_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0238_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0239_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0240_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0241_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0242_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0243_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0244_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0245_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0246_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0247_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0248_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0249_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0250_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0251_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0252_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0253_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0254_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0255_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0256_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0257_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0258_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0259_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0260_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0261_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0262_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0263_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0264_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0265_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0266_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0267_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0268_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0269_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0270_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0271_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0272_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0273_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0274_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0275_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0276_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0277_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0278_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0279_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0280_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0281_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0282_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0283_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0284_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0285_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0286_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0287_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0288_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0289_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0290_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0291_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0292_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0293_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0294_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0295_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0296_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0297_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0298_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0299_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0300_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0301_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0302_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0303_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0304_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0305_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0306_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0307_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0308_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0309_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0310_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0311_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0312_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0313_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0314_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0315_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0316_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0317_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0318_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0319_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0320_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0321_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0322_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0323_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0324_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0325_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0326_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0327_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0328_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0329_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0330_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0331_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0332_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0333_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0334_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0335_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0336_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0337_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0338_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0339_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0340_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0341_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0342_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0343_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0344_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0345_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0346_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0347_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0348_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0349_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0350_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0351_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0352_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0353_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0354_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0355_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0356_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0357_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0358_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0359_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0360_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0361_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0362_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0363_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0364_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0365_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0366_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0367_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0368_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0369_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0370_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0371_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0372_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0373_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0374_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0375_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0376_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0377_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0378_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0379_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0380_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0381_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0382_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0383_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0384_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0385_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0386_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0387_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0388_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0389_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0390_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0391_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0392_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0393_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0394_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0395_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0396_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0397_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0398_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0399_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0400_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0401_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0402_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0403_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0404_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0405_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0406_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0407_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0408_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0409_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0410_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0411_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0412_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0413_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0414_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0415_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0416_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0417_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0418_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0419_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0420_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0421_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0422_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0423_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0424_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0425_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0426_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0427_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0428_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0429_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0430_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0431_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0432_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0433_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0434_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0435_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0436_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0437_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0438_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0439_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0440_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0441_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0442_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0443_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0444_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0445_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0446_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0447_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0448_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0449_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0450_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0451_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0452_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0453_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0454_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0455_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0456_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0457_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0458_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0459_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0460_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0461_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0462_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0463_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0464_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0465_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0466_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0467_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0468_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0469_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0470_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0471_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0472_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0473_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0474_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0475_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0476_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0477_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0478_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0479_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0480_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0481_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0482_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0483_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0484_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0485_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0486_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0487_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0488_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0489_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0490_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0491_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0492_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0493_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0494_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0495_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0496_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0497_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0498_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0499_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0500_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0501_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0502_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0503_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0504_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0505_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0506_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0507_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0508_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0509_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0510_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0511_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0512_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0513_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0514_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0515_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0516_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0517_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0518_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0519_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0520_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0521_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0522_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0523_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0524_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0525_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0526_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0527_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0528_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0529_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0530_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0531_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0532_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0533_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0534_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0535_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0536_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0537_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0538_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0539_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0540_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0541_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0542_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0543_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0544_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0545_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0546_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0547_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0548_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0549_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0550_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0551_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0552_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0553_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0554_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0555_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0556_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0557_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0558_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0559_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0560_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0561_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0562_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0563_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0564_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0565_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0566_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0567_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0568_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0569_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0570_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0571_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0572_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0573_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0574_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0575_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0576_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0577_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0578_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0579_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0580_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0581_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0582_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0583_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0584_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0585_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0586_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0587_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0588_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0589_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0590_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0591_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0592_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0593_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0594_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0595_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0596_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0597_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0598_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0599_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0600_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0601_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0602_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0603_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0604_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0605_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0606_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0607_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0608_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0609_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0610_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0611_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0612_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0613_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0614_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0615_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0616_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0617_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0618_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0619_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0620_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0621_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0622_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0623_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0624_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0625_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0626_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0627_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0628_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0629_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0630_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0631_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0632_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0633_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0634_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0635_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0636_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0637_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0638_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0639_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0640_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0641_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0642_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0643_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0644_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0645_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0646_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0647_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0648_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0649_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0650_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0651_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0652_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0653_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0654_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0655_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0656_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0657_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0658_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0659_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0660_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0661_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0662_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0663_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0664_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0665_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0666_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0667_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0668_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0669_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0670_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0671_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0672_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0673_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0674_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0675_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0676_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0677_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0678_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0679_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0680_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0681_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0682_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0683_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0684_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0685_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0686_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0687_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0688_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0689_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0690_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0691_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0692_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0693_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0694_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0695_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0696_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0697_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0698_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0699_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0700_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0701_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0702_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0703_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0704_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0705_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0706_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0707_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0708_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0709_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0710_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0711_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0712_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0713_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0714_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0715_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0716_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0717_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0718_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0719_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0720_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0721_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0722_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0723_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0724_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0725_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0726_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0727_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0728_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0729_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0730_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0731_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0732_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0733_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0734_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0735_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0736_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0737_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0738_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0739_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0740_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0741_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0742_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0743_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0744_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0745_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0746_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0747_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0748_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0749_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0750_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0751_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0752_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0753_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0754_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0755_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0756_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0757_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0758_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0759_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0760_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0761_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0762_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0763_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0764_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0765_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0766_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0767_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0768_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0769_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0770_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0771_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0772_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0773_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0774_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0775_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0776_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0777_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0778_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0779_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0780_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0781_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0782_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0783_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0784_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0785_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0786_ ;
 wire \u_usb_host.u_core.u_fifo_tx._0787_ ;
 wire \u_usb_host.u_core.u_fifo_tx.count[0] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[1] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[2] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[3] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[4] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[5] ;
 wire \u_usb_host.u_core.u_fifo_tx.count[6] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[0] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[1] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[2] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[3] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[4] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[5] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[6] ;
 wire \u_usb_host.u_core.u_fifo_tx.data_i[7] ;
 wire \u_usb_host.u_core.u_fifo_tx.flush_i ;
 wire \u_usb_host.u_core.u_fifo_tx.push_i ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[0][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[10][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[11][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[12][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[13][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[14][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[15][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[16][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[17][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[18][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[19][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[1][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[20][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[21][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[22][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[23][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[24][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[25][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[26][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[27][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[28][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[29][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[2][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[30][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[31][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[32][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[33][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[34][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[35][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[36][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[37][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[38][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[39][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[3][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[40][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[41][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[42][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[43][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[44][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[45][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[46][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[47][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[48][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[49][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[4][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[50][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[51][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[52][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[53][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[54][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[55][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[56][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[57][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[58][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[59][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[5][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[60][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[61][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[62][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[63][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[6][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[7][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[8][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][0] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][1] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][2] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][3] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][4] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][5] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][6] ;
 wire \u_usb_host.u_core.u_fifo_tx.ram[9][7] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[0] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[1] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[3] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ;
 wire \u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ;
 wire \u_usb_host.u_core.u_sie._000_ ;
 wire \u_usb_host.u_core.u_sie._001_ ;
 wire \u_usb_host.u_core.u_sie._002_ ;
 wire \u_usb_host.u_core.u_sie._003_ ;
 wire \u_usb_host.u_core.u_sie._004_ ;
 wire \u_usb_host.u_core.u_sie._005_ ;
 wire \u_usb_host.u_core.u_sie._006_ ;
 wire \u_usb_host.u_core.u_sie._007_ ;
 wire \u_usb_host.u_core.u_sie._008_ ;
 wire \u_usb_host.u_core.u_sie._009_ ;
 wire \u_usb_host.u_core.u_sie._010_ ;
 wire \u_usb_host.u_core.u_sie._011_ ;
 wire \u_usb_host.u_core.u_sie._012_ ;
 wire \u_usb_host.u_core.u_sie._013_ ;
 wire \u_usb_host.u_core.u_sie._014_ ;
 wire \u_usb_host.u_core.u_sie._015_ ;
 wire \u_usb_host.u_core.u_sie._016_ ;
 wire \u_usb_host.u_core.u_sie._017_ ;
 wire \u_usb_host.u_core.u_sie._018_ ;
 wire \u_usb_host.u_core.u_sie._019_ ;
 wire \u_usb_host.u_core.u_sie._020_ ;
 wire \u_usb_host.u_core.u_sie._021_ ;
 wire \u_usb_host.u_core.u_sie._022_ ;
 wire \u_usb_host.u_core.u_sie._023_ ;
 wire \u_usb_host.u_core.u_sie._024_ ;
 wire \u_usb_host.u_core.u_sie._025_ ;
 wire \u_usb_host.u_core.u_sie._026_ ;
 wire \u_usb_host.u_core.u_sie._027_ ;
 wire \u_usb_host.u_core.u_sie._028_ ;
 wire \u_usb_host.u_core.u_sie._029_ ;
 wire \u_usb_host.u_core.u_sie._030_ ;
 wire \u_usb_host.u_core.u_sie._031_ ;
 wire \u_usb_host.u_core.u_sie._032_ ;
 wire \u_usb_host.u_core.u_sie._033_ ;
 wire \u_usb_host.u_core.u_sie._034_ ;
 wire \u_usb_host.u_core.u_sie._035_ ;
 wire \u_usb_host.u_core.u_sie._036_ ;
 wire \u_usb_host.u_core.u_sie._037_ ;
 wire \u_usb_host.u_core.u_sie._038_ ;
 wire \u_usb_host.u_core.u_sie._039_ ;
 wire \u_usb_host.u_core.u_sie._040_ ;
 wire \u_usb_host.u_core.u_sie._041_ ;
 wire \u_usb_host.u_core.u_sie._042_ ;
 wire \u_usb_host.u_core.u_sie._043_ ;
 wire \u_usb_host.u_core.u_sie._044_ ;
 wire \u_usb_host.u_core.u_sie._045_ ;
 wire \u_usb_host.u_core.u_sie._046_ ;
 wire \u_usb_host.u_core.u_sie._047_ ;
 wire \u_usb_host.u_core.u_sie._048_ ;
 wire \u_usb_host.u_core.u_sie._049_ ;
 wire \u_usb_host.u_core.u_sie._050_ ;
 wire \u_usb_host.u_core.u_sie._051_ ;
 wire \u_usb_host.u_core.u_sie._052_ ;
 wire \u_usb_host.u_core.u_sie._053_ ;
 wire \u_usb_host.u_core.u_sie._054_ ;
 wire \u_usb_host.u_core.u_sie._055_ ;
 wire \u_usb_host.u_core.u_sie._056_ ;
 wire \u_usb_host.u_core.u_sie._057_ ;
 wire \u_usb_host.u_core.u_sie._058_ ;
 wire \u_usb_host.u_core.u_sie._059_ ;
 wire \u_usb_host.u_core.u_sie._060_ ;
 wire \u_usb_host.u_core.u_sie._061_ ;
 wire \u_usb_host.u_core.u_sie._062_ ;
 wire \u_usb_host.u_core.u_sie._063_ ;
 wire \u_usb_host.u_core.u_sie._064_ ;
 wire \u_usb_host.u_core.u_sie._065_ ;
 wire \u_usb_host.u_core.u_sie._066_ ;
 wire \u_usb_host.u_core.u_sie._067_ ;
 wire \u_usb_host.u_core.u_sie._068_ ;
 wire \u_usb_host.u_core.u_sie._069_ ;
 wire \u_usb_host.u_core.u_sie._070_ ;
 wire \u_usb_host.u_core.u_sie._071_ ;
 wire \u_usb_host.u_core.u_sie._072_ ;
 wire \u_usb_host.u_core.u_sie._073_ ;
 wire \u_usb_host.u_core.u_sie._074_ ;
 wire \u_usb_host.u_core.u_sie._075_ ;
 wire \u_usb_host.u_core.u_sie._076_ ;
 wire \u_usb_host.u_core.u_sie._077_ ;
 wire \u_usb_host.u_core.u_sie._078_ ;
 wire \u_usb_host.u_core.u_sie._079_ ;
 wire \u_usb_host.u_core.u_sie._080_ ;
 wire \u_usb_host.u_core.u_sie._081_ ;
 wire \u_usb_host.u_core.u_sie._082_ ;
 wire \u_usb_host.u_core.u_sie._083_ ;
 wire \u_usb_host.u_core.u_sie._084_ ;
 wire \u_usb_host.u_core.u_sie._085_ ;
 wire \u_usb_host.u_core.u_sie._086_ ;
 wire \u_usb_host.u_core.u_sie._087_ ;
 wire \u_usb_host.u_core.u_sie._088_ ;
 wire \u_usb_host.u_core.u_sie._089_ ;
 wire \u_usb_host.u_core.u_sie._090_ ;
 wire \u_usb_host.u_core.u_sie._091_ ;
 wire \u_usb_host.u_core.u_sie._092_ ;
 wire \u_usb_host.u_core.u_sie._093_ ;
 wire \u_usb_host.u_core.u_sie._094_ ;
 wire \u_usb_host.u_core.u_sie._095_ ;
 wire \u_usb_host.u_core.u_sie._096_ ;
 wire \u_usb_host.u_core.u_sie._097_ ;
 wire \u_usb_host.u_core.u_sie._098_ ;
 wire \u_usb_host.u_core.u_sie._099_ ;
 wire \u_usb_host.u_core.u_sie._100_ ;
 wire \u_usb_host.u_core.u_sie._101_ ;
 wire \u_usb_host.u_core.u_sie._102_ ;
 wire \u_usb_host.u_core.u_sie._103_ ;
 wire \u_usb_host.u_core.u_sie._104_ ;
 wire \u_usb_host.u_core.u_sie._105_ ;
 wire \u_usb_host.u_core.u_sie._106_ ;
 wire \u_usb_host.u_core.u_sie._107_ ;
 wire \u_usb_host.u_core.u_sie._108_ ;
 wire \u_usb_host.u_core.u_sie._109_ ;
 wire \u_usb_host.u_core.u_sie._110_ ;
 wire \u_usb_host.u_core.u_sie._111_ ;
 wire \u_usb_host.u_core.u_sie._112_ ;
 wire \u_usb_host.u_core.u_sie._113_ ;
 wire \u_usb_host.u_core.u_sie._114_ ;
 wire \u_usb_host.u_core.u_sie._115_ ;
 wire \u_usb_host.u_core.u_sie._116_ ;
 wire \u_usb_host.u_core.u_sie._117_ ;
 wire \u_usb_host.u_core.u_sie._118_ ;
 wire \u_usb_host.u_core.u_sie._119_ ;
 wire \u_usb_host.u_core.u_sie._120_ ;
 wire \u_usb_host.u_core.u_sie._121_ ;
 wire \u_usb_host.u_core.u_sie._122_ ;
 wire \u_usb_host.u_core.u_sie._123_ ;
 wire \u_usb_host.u_core.u_sie._124_ ;
 wire \u_usb_host.u_core.u_sie._125_ ;
 wire \u_usb_host.u_core.u_sie._126_ ;
 wire \u_usb_host.u_core.u_sie._127_ ;
 wire \u_usb_host.u_core.u_sie._128_ ;
 wire \u_usb_host.u_core.u_sie._129_ ;
 wire \u_usb_host.u_core.u_sie._130_ ;
 wire \u_usb_host.u_core.u_sie._131_ ;
 wire \u_usb_host.u_core.u_sie._132_ ;
 wire \u_usb_host.u_core.u_sie._133_ ;
 wire \u_usb_host.u_core.u_sie._134_ ;
 wire \u_usb_host.u_core.u_sie._135_ ;
 wire \u_usb_host.u_core.u_sie._136_ ;
 wire \u_usb_host.u_core.u_sie._137_ ;
 wire \u_usb_host.u_core.u_sie._138_ ;
 wire \u_usb_host.u_core.u_sie._139_ ;
 wire \u_usb_host.u_core.u_sie._140_ ;
 wire \u_usb_host.u_core.u_sie._141_ ;
 wire \u_usb_host.u_core.u_sie._142_ ;
 wire \u_usb_host.u_core.u_sie._143_ ;
 wire \u_usb_host.u_core.u_sie._144_ ;
 wire \u_usb_host.u_core.u_sie._145_ ;
 wire \u_usb_host.u_core.u_sie._146_ ;
 wire \u_usb_host.u_core.u_sie._147_ ;
 wire \u_usb_host.u_core.u_sie._148_ ;
 wire \u_usb_host.u_core.u_sie._149_ ;
 wire \u_usb_host.u_core.u_sie._150_ ;
 wire \u_usb_host.u_core.u_sie._151_ ;
 wire \u_usb_host.u_core.u_sie._152_ ;
 wire \u_usb_host.u_core.u_sie._153_ ;
 wire \u_usb_host.u_core.u_sie._154_ ;
 wire \u_usb_host.u_core.u_sie._155_ ;
 wire \u_usb_host.u_core.u_sie._156_ ;
 wire \u_usb_host.u_core.u_sie._157_ ;
 wire \u_usb_host.u_core.u_sie._158_ ;
 wire \u_usb_host.u_core.u_sie._159_ ;
 wire \u_usb_host.u_core.u_sie._160_ ;
 wire \u_usb_host.u_core.u_sie._161_ ;
 wire \u_usb_host.u_core.u_sie._162_ ;
 wire \u_usb_host.u_core.u_sie._163_ ;
 wire \u_usb_host.u_core.u_sie._164_ ;
 wire \u_usb_host.u_core.u_sie._165_ ;
 wire \u_usb_host.u_core.u_sie._166_ ;
 wire \u_usb_host.u_core.u_sie._167_ ;
 wire \u_usb_host.u_core.u_sie._168_ ;
 wire \u_usb_host.u_core.u_sie._169_ ;
 wire \u_usb_host.u_core.u_sie._170_ ;
 wire \u_usb_host.u_core.u_sie._171_ ;
 wire \u_usb_host.u_core.u_sie._172_ ;
 wire \u_usb_host.u_core.u_sie._173_ ;
 wire \u_usb_host.u_core.u_sie._174_ ;
 wire \u_usb_host.u_core.u_sie._175_ ;
 wire \u_usb_host.u_core.u_sie._176_ ;
 wire \u_usb_host.u_core.u_sie._177_ ;
 wire \u_usb_host.u_core.u_sie._178_ ;
 wire \u_usb_host.u_core.u_sie._179_ ;
 wire \u_usb_host.u_core.u_sie._180_ ;
 wire \u_usb_host.u_core.u_sie._181_ ;
 wire \u_usb_host.u_core.u_sie._182_ ;
 wire \u_usb_host.u_core.u_sie._183_ ;
 wire \u_usb_host.u_core.u_sie._184_ ;
 wire \u_usb_host.u_core.u_sie._185_ ;
 wire \u_usb_host.u_core.u_sie._186_ ;
 wire \u_usb_host.u_core.u_sie._187_ ;
 wire \u_usb_host.u_core.u_sie._188_ ;
 wire \u_usb_host.u_core.u_sie._189_ ;
 wire \u_usb_host.u_core.u_sie._190_ ;
 wire \u_usb_host.u_core.u_sie._191_ ;
 wire \u_usb_host.u_core.u_sie._192_ ;
 wire \u_usb_host.u_core.u_sie._193_ ;
 wire \u_usb_host.u_core.u_sie._194_ ;
 wire \u_usb_host.u_core.u_sie._195_ ;
 wire \u_usb_host.u_core.u_sie._196_ ;
 wire \u_usb_host.u_core.u_sie._197_ ;
 wire \u_usb_host.u_core.u_sie._198_ ;
 wire \u_usb_host.u_core.u_sie._199_ ;
 wire \u_usb_host.u_core.u_sie._200_ ;
 wire \u_usb_host.u_core.u_sie._201_ ;
 wire \u_usb_host.u_core.u_sie._202_ ;
 wire \u_usb_host.u_core.u_sie._203_ ;
 wire \u_usb_host.u_core.u_sie._204_ ;
 wire \u_usb_host.u_core.u_sie._205_ ;
 wire \u_usb_host.u_core.u_sie._206_ ;
 wire \u_usb_host.u_core.u_sie._207_ ;
 wire \u_usb_host.u_core.u_sie._208_ ;
 wire \u_usb_host.u_core.u_sie._209_ ;
 wire \u_usb_host.u_core.u_sie._210_ ;
 wire \u_usb_host.u_core.u_sie._211_ ;
 wire \u_usb_host.u_core.u_sie._212_ ;
 wire \u_usb_host.u_core.u_sie._213_ ;
 wire \u_usb_host.u_core.u_sie._214_ ;
 wire \u_usb_host.u_core.u_sie._215_ ;
 wire \u_usb_host.u_core.u_sie._216_ ;
 wire \u_usb_host.u_core.u_sie._217_ ;
 wire \u_usb_host.u_core.u_sie._218_ ;
 wire \u_usb_host.u_core.u_sie._219_ ;
 wire \u_usb_host.u_core.u_sie._220_ ;
 wire \u_usb_host.u_core.u_sie._221_ ;
 wire \u_usb_host.u_core.u_sie._222_ ;
 wire \u_usb_host.u_core.u_sie._223_ ;
 wire \u_usb_host.u_core.u_sie._224_ ;
 wire \u_usb_host.u_core.u_sie._225_ ;
 wire \u_usb_host.u_core.u_sie._226_ ;
 wire \u_usb_host.u_core.u_sie._227_ ;
 wire \u_usb_host.u_core.u_sie._228_ ;
 wire \u_usb_host.u_core.u_sie._229_ ;
 wire \u_usb_host.u_core.u_sie._230_ ;
 wire \u_usb_host.u_core.u_sie._231_ ;
 wire \u_usb_host.u_core.u_sie._232_ ;
 wire \u_usb_host.u_core.u_sie._233_ ;
 wire \u_usb_host.u_core.u_sie._234_ ;
 wire \u_usb_host.u_core.u_sie._235_ ;
 wire \u_usb_host.u_core.u_sie._236_ ;
 wire \u_usb_host.u_core.u_sie._237_ ;
 wire \u_usb_host.u_core.u_sie._238_ ;
 wire \u_usb_host.u_core.u_sie._239_ ;
 wire \u_usb_host.u_core.u_sie._240_ ;
 wire \u_usb_host.u_core.u_sie._241_ ;
 wire \u_usb_host.u_core.u_sie._242_ ;
 wire \u_usb_host.u_core.u_sie._243_ ;
 wire \u_usb_host.u_core.u_sie._244_ ;
 wire \u_usb_host.u_core.u_sie._245_ ;
 wire \u_usb_host.u_core.u_sie._246_ ;
 wire \u_usb_host.u_core.u_sie._247_ ;
 wire \u_usb_host.u_core.u_sie._248_ ;
 wire \u_usb_host.u_core.u_sie._249_ ;
 wire \u_usb_host.u_core.u_sie._250_ ;
 wire \u_usb_host.u_core.u_sie._251_ ;
 wire \u_usb_host.u_core.u_sie._252_ ;
 wire \u_usb_host.u_core.u_sie._253_ ;
 wire \u_usb_host.u_core.u_sie._254_ ;
 wire \u_usb_host.u_core.u_sie._255_ ;
 wire \u_usb_host.u_core.u_sie._256_ ;
 wire \u_usb_host.u_core.u_sie._257_ ;
 wire \u_usb_host.u_core.u_sie._258_ ;
 wire \u_usb_host.u_core.u_sie._259_ ;
 wire \u_usb_host.u_core.u_sie._260_ ;
 wire \u_usb_host.u_core.u_sie._261_ ;
 wire \u_usb_host.u_core.u_sie._262_ ;
 wire \u_usb_host.u_core.u_sie._263_ ;
 wire \u_usb_host.u_core.u_sie._264_ ;
 wire \u_usb_host.u_core.u_sie._265_ ;
 wire \u_usb_host.u_core.u_sie._266_ ;
 wire \u_usb_host.u_core.u_sie._267_ ;
 wire \u_usb_host.u_core.u_sie._268_ ;
 wire \u_usb_host.u_core.u_sie._269_ ;
 wire \u_usb_host.u_core.u_sie._270_ ;
 wire \u_usb_host.u_core.u_sie._271_ ;
 wire \u_usb_host.u_core.u_sie._272_ ;
 wire \u_usb_host.u_core.u_sie._273_ ;
 wire \u_usb_host.u_core.u_sie._274_ ;
 wire \u_usb_host.u_core.u_sie._275_ ;
 wire \u_usb_host.u_core.u_sie._276_ ;
 wire \u_usb_host.u_core.u_sie._277_ ;
 wire \u_usb_host.u_core.u_sie._278_ ;
 wire \u_usb_host.u_core.u_sie._279_ ;
 wire \u_usb_host.u_core.u_sie._280_ ;
 wire \u_usb_host.u_core.u_sie._281_ ;
 wire \u_usb_host.u_core.u_sie._282_ ;
 wire \u_usb_host.u_core.u_sie._283_ ;
 wire \u_usb_host.u_core.u_sie._284_ ;
 wire \u_usb_host.u_core.u_sie._285_ ;
 wire \u_usb_host.u_core.u_sie._286_ ;
 wire \u_usb_host.u_core.u_sie._287_ ;
 wire \u_usb_host.u_core.u_sie._288_ ;
 wire \u_usb_host.u_core.u_sie._289_ ;
 wire \u_usb_host.u_core.u_sie._290_ ;
 wire \u_usb_host.u_core.u_sie._291_ ;
 wire \u_usb_host.u_core.u_sie._292_ ;
 wire \u_usb_host.u_core.u_sie._293_ ;
 wire \u_usb_host.u_core.u_sie._294_ ;
 wire \u_usb_host.u_core.u_sie._295_ ;
 wire \u_usb_host.u_core.u_sie._296_ ;
 wire \u_usb_host.u_core.u_sie._297_ ;
 wire \u_usb_host.u_core.u_sie._298_ ;
 wire \u_usb_host.u_core.u_sie._299_ ;
 wire \u_usb_host.u_core.u_sie._300_ ;
 wire \u_usb_host.u_core.u_sie._301_ ;
 wire \u_usb_host.u_core.u_sie._302_ ;
 wire \u_usb_host.u_core.u_sie._303_ ;
 wire \u_usb_host.u_core.u_sie._304_ ;
 wire \u_usb_host.u_core.u_sie._305_ ;
 wire \u_usb_host.u_core.u_sie._306_ ;
 wire \u_usb_host.u_core.u_sie._307_ ;
 wire \u_usb_host.u_core.u_sie._308_ ;
 wire \u_usb_host.u_core.u_sie._309_ ;
 wire \u_usb_host.u_core.u_sie._310_ ;
 wire \u_usb_host.u_core.u_sie._311_ ;
 wire \u_usb_host.u_core.u_sie._312_ ;
 wire \u_usb_host.u_core.u_sie.crc5_out_w[0] ;
 wire \u_usb_host.u_core.u_sie.crc5_out_w[1] ;
 wire \u_usb_host.u_core.u_sie.crc5_out_w[2] ;
 wire \u_usb_host.u_core.u_sie.crc5_out_w[3] ;
 wire \u_usb_host.u_core.u_sie.crc5_out_w[4] ;
 wire \u_usb_host.u_core.u_sie.crc_byte_w ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[0] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[1] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[2] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[3] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[4] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[5] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[6] ;
 wire \u_usb_host.u_core.u_sie.crc_data_in_w[7] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[0] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[10] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[11] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[12] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[13] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[14] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[15] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[1] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[2] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[3] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[4] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[5] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[6] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[7] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[8] ;
 wire \u_usb_host.u_core.u_sie.crc_out_w[9] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[0] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[10] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[11] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[12] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[13] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[14] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[15] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[1] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[2] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[3] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[4] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[5] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[6] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[7] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[8] ;
 wire \u_usb_host.u_core.u_sie.crc_sum_q[9] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[0] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[10] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[11] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[12] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[13] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[14] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[15] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[16] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[17] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[18] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[19] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[1] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[20] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[21] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[22] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[23] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[24] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[25] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[26] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[27] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[28] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[29] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[2] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[30] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[31] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[3] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[4] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[5] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[6] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[7] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[8] ;
 wire \u_usb_host.u_core.u_sie.data_buffer_q[9] ;
 wire \u_usb_host.u_core.u_sie.data_crc_q[1] ;
 wire \u_usb_host.u_core.u_sie.data_idx_i ;
 wire \u_usb_host.u_core.u_sie.data_len_i[0] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[10] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[11] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[12] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[13] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[14] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[15] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[1] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[2] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[3] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[4] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[5] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[6] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[7] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[8] ;
 wire \u_usb_host.u_core.u_sie.data_len_i[9] ;
 wire \u_usb_host.u_core.u_sie.data_ready_w ;
 wire \u_usb_host.u_core.u_sie.data_valid_q[1] ;
 wire \u_usb_host.u_core.u_sie.data_valid_q[2] ;
 wire \u_usb_host.u_core.u_sie.data_valid_q[3] ;
 wire \u_usb_host.u_core.u_sie.in_transfer_q ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[0] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[1] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[2] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[3] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[4] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[5] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[6] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[7] ;
 wire \u_usb_host.u_core.u_sie.last_tx_time_q[8] ;
 wire \u_usb_host.u_core.u_sie.next_state_r[0] ;
 wire \u_usb_host.u_core.u_sie.next_state_r[1] ;
 wire \u_usb_host.u_core.u_sie.next_state_r[2] ;
 wire \u_usb_host.u_core.u_sie.next_state_r[3] ;
 wire \u_usb_host.u_core.u_sie.rx_active_q[0] ;
 wire \u_usb_host.u_core.u_sie.rx_active_q[1] ;
 wire \u_usb_host.u_core.u_sie.rx_active_q[2] ;
 wire \u_usb_host.u_core.u_sie.rx_active_q[3] ;
 wire \u_usb_host.u_core.u_sie.se0_detect_q ;
 wire \u_usb_host.u_core.u_sie.se0_detect_w ;
 wire \u_usb_host.u_core.u_sie.send_ack_q ;
 wire \u_usb_host.u_core.u_sie.send_data1_q ;
 wire \u_usb_host.u_core.u_sie.send_sof_q ;
 wire \u_usb_host.u_core.u_sie.shift_en_w ;
 wire \u_usb_host.u_core.u_sie.state_q[0] ;
 wire \u_usb_host.u_core.u_sie.state_q[1] ;
 wire \u_usb_host.u_core.u_sie.state_q[2] ;
 wire \u_usb_host.u_core.u_sie.state_q[3] ;
 wire \u_usb_host.u_core.u_sie.token_q[0] ;
 wire \u_usb_host.u_core.u_sie.token_q[10] ;
 wire \u_usb_host.u_core.u_sie.token_q[11] ;
 wire \u_usb_host.u_core.u_sie.token_q[12] ;
 wire \u_usb_host.u_core.u_sie.token_q[13] ;
 wire \u_usb_host.u_core.u_sie.token_q[14] ;
 wire \u_usb_host.u_core.u_sie.token_q[15] ;
 wire \u_usb_host.u_core.u_sie.token_q[1] ;
 wire \u_usb_host.u_core.u_sie.token_q[2] ;
 wire \u_usb_host.u_core.u_sie.token_q[3] ;
 wire \u_usb_host.u_core.u_sie.token_q[4] ;
 wire \u_usb_host.u_core.u_sie.token_q[5] ;
 wire \u_usb_host.u_core.u_sie.token_q[6] ;
 wire \u_usb_host.u_core.u_sie.token_q[7] ;
 wire \u_usb_host.u_core.u_sie.token_q[8] ;
 wire \u_usb_host.u_core.u_sie.token_q[9] ;
 wire \u_usb_host.u_core.u_sie.tx_ifs_q[0] ;
 wire \u_usb_host.u_core.u_sie.tx_ifs_q[1] ;
 wire \u_usb_host.u_core.u_sie.tx_ifs_q[2] ;
 wire \u_usb_host.u_core.u_sie.tx_ifs_q[3] ;
 wire \u_usb_host.u_core.u_sie.u_crc16._00_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._01_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._02_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._03_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._04_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._05_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._06_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._07_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._08_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._09_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._10_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._11_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._12_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._13_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._14_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._15_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._16_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._17_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._18_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._19_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._20_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._21_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._22_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._23_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._24_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._25_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._26_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._27_ ;
 wire \u_usb_host.u_core.u_sie.u_crc16._28_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._00_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._01_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._02_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._03_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._04_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._05_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._06_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._07_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._08_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._09_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._10_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._11_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._12_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._13_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._14_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._15_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._16_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._17_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._18_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._19_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._20_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._21_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._22_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._23_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._24_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._25_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._26_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._27_ ;
 wire \u_usb_host.u_core.u_sie.u_crc5._28_ ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[2] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[3] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[4] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[5] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[6] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_i[7] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[2] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[3] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[4] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[5] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[6] ;
 wire \u_usb_host.u_core.u_sie.utmi_data_o[7] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_i[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_i[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_q[0] ;
 wire \u_usb_host.u_core.u_sie.utmi_linestate_q[1] ;
 wire \u_usb_host.u_core.u_sie.utmi_rxactive_i ;
 wire \u_usb_host.u_core.u_sie.utmi_rxvalid_i ;
 wire \u_usb_host.u_core.u_sie.utmi_txready_i ;
 wire \u_usb_host.u_core.u_sie.utmi_txvalid_o ;
 wire \u_usb_host.u_core.u_sie.wait_eop_q ;
 wire \u_usb_host.u_core.u_sie.wait_resp_q ;
 wire \u_usb_host.u_core.usb_ctrl_enable_sof_out_w ;
 wire \u_usb_host.u_core.usb_ctrl_wr_q ;
 wire \u_usb_host.u_core.usb_err_q ;
 wire \u_usb_host.u_core.usb_irq_ack_device_detect_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_done_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_err_out_w ;
 wire \u_usb_host.u_core.usb_irq_ack_sof_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_device_detect_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_done_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_err_out_w ;
 wire \u_usb_host.u_core.usb_irq_mask_sof_out_w ;
 wire \u_usb_host.u_core.usb_rx_stat_start_pend_in_w ;
 wire \u_usb_host.u_core.usb_xfer_token_ack_out_w ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ;
 wire \u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_in_out_w ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ;
 wire \u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ;
 wire \u_usb_host.u_core.utmi_dmpulldown_o ;
 wire \u_usb_host.u_core.utmi_dppulldown_o ;
 wire \u_usb_host.u_core.utmi_op_mode_o[0] ;
 wire \u_usb_host.u_core.utmi_op_mode_o[1] ;
 wire \u_usb_host.u_core.utmi_rxerror_i ;
 wire \u_usb_host.u_core.utmi_termselect_o ;
 wire \u_usb_host.u_core.utmi_xcvrselect_o[0] ;
 wire \u_usb_host.u_core.utmi_xcvrselect_o[1] ;
 wire \u_usb_host.u_phy._000_ ;
 wire \u_usb_host.u_phy._001_ ;
 wire \u_usb_host.u_phy._002_ ;
 wire \u_usb_host.u_phy._003_ ;
 wire \u_usb_host.u_phy._004_ ;
 wire \u_usb_host.u_phy._005_ ;
 wire \u_usb_host.u_phy._006_ ;
 wire \u_usb_host.u_phy._007_ ;
 wire \u_usb_host.u_phy._008_ ;
 wire \u_usb_host.u_phy._009_ ;
 wire \u_usb_host.u_phy._010_ ;
 wire \u_usb_host.u_phy._011_ ;
 wire \u_usb_host.u_phy._012_ ;
 wire \u_usb_host.u_phy._013_ ;
 wire \u_usb_host.u_phy._014_ ;
 wire \u_usb_host.u_phy._015_ ;
 wire \u_usb_host.u_phy._016_ ;
 wire \u_usb_host.u_phy._017_ ;
 wire \u_usb_host.u_phy._018_ ;
 wire \u_usb_host.u_phy._019_ ;
 wire \u_usb_host.u_phy._020_ ;
 wire \u_usb_host.u_phy._021_ ;
 wire \u_usb_host.u_phy._022_ ;
 wire \u_usb_host.u_phy._030_ ;
 wire \u_usb_host.u_phy._031_ ;
 wire \u_usb_host.u_phy._032_ ;
 wire \u_usb_host.u_phy._033_ ;
 wire \u_usb_host.u_phy._034_ ;
 wire \u_usb_host.u_phy._036_ ;
 wire \u_usb_host.u_phy._037_ ;
 wire \u_usb_host.u_phy._038_ ;
 wire \u_usb_host.u_phy._039_ ;
 wire \u_usb_host.u_phy._040_ ;
 wire \u_usb_host.u_phy._041_ ;
 wire \u_usb_host.u_phy._042_ ;
 wire \u_usb_host.u_phy._043_ ;
 wire \u_usb_host.u_phy._045_ ;
 wire \u_usb_host.u_phy._046_ ;
 wire \u_usb_host.u_phy._047_ ;
 wire \u_usb_host.u_phy._048_ ;
 wire \u_usb_host.u_phy._049_ ;
 wire \u_usb_host.u_phy._050_ ;
 wire \u_usb_host.u_phy._051_ ;
 wire \u_usb_host.u_phy._052_ ;
 wire \u_usb_host.u_phy._053_ ;
 wire \u_usb_host.u_phy._054_ ;
 wire \u_usb_host.u_phy._055_ ;
 wire \u_usb_host.u_phy._056_ ;
 wire \u_usb_host.u_phy._057_ ;
 wire \u_usb_host.u_phy._058_ ;
 wire \u_usb_host.u_phy._059_ ;
 wire \u_usb_host.u_phy._060_ ;
 wire \u_usb_host.u_phy._061_ ;
 wire \u_usb_host.u_phy._062_ ;
 wire \u_usb_host.u_phy._063_ ;
 wire \u_usb_host.u_phy._064_ ;
 wire \u_usb_host.u_phy._065_ ;
 wire \u_usb_host.u_phy._066_ ;
 wire \u_usb_host.u_phy._067_ ;
 wire \u_usb_host.u_phy._068_ ;
 wire \u_usb_host.u_phy._069_ ;
 wire \u_usb_host.u_phy._070_ ;
 wire \u_usb_host.u_phy._071_ ;
 wire \u_usb_host.u_phy._072_ ;
 wire \u_usb_host.u_phy._073_ ;
 wire \u_usb_host.u_phy._074_ ;
 wire \u_usb_host.u_phy._075_ ;
 wire \u_usb_host.u_phy._076_ ;
 wire \u_usb_host.u_phy._077_ ;
 wire \u_usb_host.u_phy._078_ ;
 wire \u_usb_host.u_phy._079_ ;
 wire \u_usb_host.u_phy._080_ ;
 wire \u_usb_host.u_phy._081_ ;
 wire \u_usb_host.u_phy._082_ ;
 wire \u_usb_host.u_phy._083_ ;
 wire \u_usb_host.u_phy._084_ ;
 wire \u_usb_host.u_phy._085_ ;
 wire \u_usb_host.u_phy._086_ ;
 wire \u_usb_host.u_phy._087_ ;
 wire \u_usb_host.u_phy._088_ ;
 wire \u_usb_host.u_phy._089_ ;
 wire \u_usb_host.u_phy._090_ ;
 wire \u_usb_host.u_phy._091_ ;
 wire \u_usb_host.u_phy._092_ ;
 wire \u_usb_host.u_phy._093_ ;
 wire \u_usb_host.u_phy._094_ ;
 wire \u_usb_host.u_phy._095_ ;
 wire \u_usb_host.u_phy._096_ ;
 wire \u_usb_host.u_phy._097_ ;
 wire \u_usb_host.u_phy._098_ ;
 wire \u_usb_host.u_phy._099_ ;
 wire \u_usb_host.u_phy._100_ ;
 wire \u_usb_host.u_phy._101_ ;
 wire \u_usb_host.u_phy._102_ ;
 wire \u_usb_host.u_phy._103_ ;
 wire \u_usb_host.u_phy._104_ ;
 wire \u_usb_host.u_phy._105_ ;
 wire \u_usb_host.u_phy._106_ ;
 wire \u_usb_host.u_phy._107_ ;
 wire \u_usb_host.u_phy._108_ ;
 wire \u_usb_host.u_phy._109_ ;
 wire \u_usb_host.u_phy._110_ ;
 wire \u_usb_host.u_phy._113_ ;
 wire \u_usb_host.u_phy._114_ ;
 wire \u_usb_host.u_phy._115_ ;
 wire \u_usb_host.u_phy._116_ ;
 wire \u_usb_host.u_phy._117_ ;
 wire \u_usb_host.u_phy._118_ ;
 wire \u_usb_host.u_phy._119_ ;
 wire \u_usb_host.u_phy._120_ ;
 wire \u_usb_host.u_phy._121_ ;
 wire \u_usb_host.u_phy._122_ ;
 wire \u_usb_host.u_phy._123_ ;
 wire \u_usb_host.u_phy._124_ ;
 wire \u_usb_host.u_phy._125_ ;
 wire \u_usb_host.u_phy._126_ ;
 wire \u_usb_host.u_phy._127_ ;
 wire \u_usb_host.u_phy._128_ ;
 wire \u_usb_host.u_phy._129_ ;
 wire \u_usb_host.u_phy._130_ ;
 wire \u_usb_host.u_phy._131_ ;
 wire \u_usb_host.u_phy._132_ ;
 wire \u_usb_host.u_phy._133_ ;
 wire \u_usb_host.u_phy._134_ ;
 wire \u_usb_host.u_phy._135_ ;
 wire \u_usb_host.u_phy._136_ ;
 wire \u_usb_host.u_phy._137_ ;
 wire \u_usb_host.u_phy._138_ ;
 wire \u_usb_host.u_phy._139_ ;
 wire \u_usb_host.u_phy._140_ ;
 wire \u_usb_host.u_phy._141_ ;
 wire \u_usb_host.u_phy._142_ ;
 wire \u_usb_host.u_phy._150_ ;
 wire \u_usb_host.u_phy._151_ ;
 wire \u_usb_host.u_phy._152_ ;
 wire \u_usb_host.u_phy._153_ ;
 wire \u_usb_host.u_phy._154_ ;
 wire \u_usb_host.u_phy._155_ ;
 wire \u_usb_host.u_phy._156_ ;
 wire \u_usb_host.u_phy._157_ ;
 wire \u_usb_host.u_phy._158_ ;
 wire \u_usb_host.u_phy._159_ ;
 wire \u_usb_host.u_phy._160_ ;
 wire \u_usb_host.u_phy._161_ ;
 wire \u_usb_host.u_phy._162_ ;
 wire \u_usb_host.u_phy._163_ ;
 wire \u_usb_host.u_phy._164_ ;
 wire \u_usb_host.u_phy._165_ ;
 wire \u_usb_host.u_phy._166_ ;
 wire \u_usb_host.u_phy._167_ ;
 wire \u_usb_host.u_phy._168_ ;
 wire \u_usb_host.u_phy._169_ ;
 wire \u_usb_host.u_phy._170_ ;
 wire \u_usb_host.u_phy._172_ ;
 wire \u_usb_host.u_phy._173_ ;
 wire \u_usb_host.u_phy._174_ ;
 wire \u_usb_host.u_phy._175_ ;
 wire \u_usb_host.u_phy._176_ ;
 wire \u_usb_host.u_phy._177_ ;
 wire \u_usb_host.u_phy._178_ ;
 wire \u_usb_host.u_phy._179_ ;
 wire \u_usb_host.u_phy._180_ ;
 wire \u_usb_host.u_phy._181_ ;
 wire \u_usb_host.u_phy._182_ ;
 wire \u_usb_host.u_phy._183_ ;
 wire \u_usb_host.u_phy.adjust_delayed_q ;
 wire \u_usb_host.u_phy.bit_count_q[0] ;
 wire \u_usb_host.u_phy.bit_count_q[1] ;
 wire \u_usb_host.u_phy.bit_count_q[2] ;
 wire \u_usb_host.u_phy.in_j_w ;
 wire \u_usb_host.u_phy.next_state_r[0] ;
 wire \u_usb_host.u_phy.next_state_r[1] ;
 wire \u_usb_host.u_phy.next_state_r[2] ;
 wire \u_usb_host.u_phy.next_state_r[3] ;
 wire \u_usb_host.u_phy.ones_count_q[0] ;
 wire \u_usb_host.u_phy.ones_count_q[1] ;
 wire \u_usb_host.u_phy.ones_count_q[2] ;
 wire \u_usb_host.u_phy.rx_dn0_q ;
 wire \u_usb_host.u_phy.rx_dn1_q ;
 wire \u_usb_host.u_phy.rx_dn_ms ;
 wire \u_usb_host.u_phy.rx_dn_q ;
 wire \u_usb_host.u_phy.rx_dp0_q ;
 wire \u_usb_host.u_phy.rx_dp1_q ;
 wire \u_usb_host.u_phy.rx_dp_ms ;
 wire \u_usb_host.u_phy.rx_dp_q ;
 wire \u_usb_host.u_phy.rxd0_q ;
 wire \u_usb_host.u_phy.rxd1_q ;
 wire \u_usb_host.u_phy.rxd_last_j_q ;
 wire \u_usb_host.u_phy.rxd_last_q ;
 wire \u_usb_host.u_phy.rxd_ms ;
 wire \u_usb_host.u_phy.rxd_q ;
 wire \u_usb_host.u_phy.sample_cnt_q[0] ;
 wire \u_usb_host.u_phy.sample_cnt_q[1] ;
 wire \u_usb_host.u_phy.sample_cnt_q[2] ;
 wire \u_usb_host.u_phy.send_eop_q ;
 wire \u_usb_host.u_phy.state_q[0] ;
 wire \u_usb_host.u_phy.state_q[1] ;
 wire \u_usb_host.u_phy.state_q[2] ;
 wire \u_usb_host.u_phy.state_q[3] ;
 wire \u_usb_host.u_phy.sync_j_detected_q ;
 wire \u_usb_host.u_phy.usb_rx_dn_i ;
 wire \u_usb_host.u_phy.usb_rx_dp_i ;
 wire \u_usb_host.u_phy.usb_rx_rcv_i ;
 wire \u_usb_host.u_phy.usb_tx_dn_o ;
 wire \u_usb_host.u_phy.usb_tx_dp_o ;
 wire \u_usb_host.u_phy.usb_tx_oen_o ;
 wire \u_usb_host.u_usb_rst.in_data_2s ;
 wire \u_usb_host.u_usb_rst.in_data_s ;
 wire \u_usb_host.u_usb_xcvr._0_ ;
 wire \u_usb_host.u_usb_xcvr._1_ ;
 wire \u_usb_host.u_wb_rst.in_data_2s ;
 wire \u_usb_host.u_wb_rst.in_data_s ;

 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_app_clk_A (.DIODE(app_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._040__A  (.DIODE(\u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_usb_clk_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_0_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_1_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_2_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_3_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_4_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_5_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_6_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_3_7_0_usb_clk_A (.DIODE(clknet_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_usb_clk_A (.DIODE(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_18_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_usb_clk_A (.DIODE(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_27_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_usb_clk_A (.DIODE(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_usb_clk_A (.DIODE(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_usb_clk_A (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_3_usb_clk_A (.DIODE(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_usb_clk_A (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_usb_clk_A (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_usb_clk_A (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_usb_clk_A (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_49_usb_clk_A (.DIODE(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_usb_clk_A (.DIODE(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_usb_clk_A (.DIODE(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_57_usb_clk_A (.DIODE(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_usb_clk_A (.DIODE(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_59_usb_clk_A (.DIODE(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_usb_clk_A (.DIODE(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_usb_clk_A (.DIODE(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout100_A (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout102_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0475_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout105_A (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout107_A (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout108_A (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout109_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout110_A (.DIODE(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout113_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout115_A (.DIODE(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout116_A (.DIODE(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout118_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout119_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout120_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout121_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout122_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout123_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout124_A (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout125_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout127_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout128_A (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout129_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout130_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout131_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout132_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout133_A (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout135_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout136_A (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout137_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout138_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout139_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout140_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout141_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout142_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout143_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout144_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout145_A (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout146_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout147_A (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout148_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout149_A (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout150_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout151_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout152_A (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout153_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout154_A (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout155_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout156_A (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout157_A (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout159_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout160_A (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout161_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout162_A (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout163_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout164_A (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout165_A (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout166_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout167_A (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout168_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout169_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout170_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout171_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout172_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout173_A (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout174_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout175_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout176_A (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout177_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout178_A (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout179_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout180_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout181_A (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout182_A (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout184_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0575_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout185_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout186_A (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout187_A (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout189_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout190_A (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout191_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0571_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout192_A (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout193_A (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout194_A (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout196_A (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout197_A (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout198_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout200_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout201_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout203_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout204_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout205_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout206_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout208_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0529_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout209_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0529_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout212_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0525_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout213_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout214_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout215_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout218_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout219_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout221_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout222_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout224_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout227_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout229_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout230_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout232_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout233_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout235_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout236_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout237_A (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout238_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout239_A (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout241_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout242_A (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout243_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0516_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout244_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout245_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout247_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout249_A (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout250_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout256_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout257_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout261_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout266_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout267_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout268_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout269_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout270_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout271_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout272_A (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout274_A (.DIODE(\u_usb_host.u_core.u_fifo_tx._0504_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout275_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0575_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout276_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0573_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout277_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0573_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout278_A (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout279_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0573_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout280_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout281_A (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout282_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0571_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout283_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout284_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout285_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout286_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout287_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout288_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout289_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout290_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout291_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout292_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout294_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout295_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0544_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout296_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout297_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout298_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0531_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout299_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0529_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout300_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0529_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout301_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0527_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout302_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout303_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0525_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout306_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout309_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout312_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout316_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout318_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout320_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout321_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout322_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout323_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout324_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout328_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout329_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout330_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout331_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout333_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout335_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout336_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout337_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout338_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout341_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout347_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout348_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout352_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout354_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout355_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout356_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout357_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout358_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0508_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout359_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout360_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout361_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout362_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout363_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0504_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout366_A (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout367_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout368_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout369_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout371_A (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout372_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout373_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout374_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout377_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout379_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout381_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout382_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout383_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout384_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout385_A (.DIODE(net386));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout386_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout388_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout389_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout390_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout391_A (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout392_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout393_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout394_A (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout395_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout397_A (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout398_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout400_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout402_A (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout403_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout404_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout405_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout406_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout408_A (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout409_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout411_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout414_A (.DIODE(net415));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout415_A (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout416_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout457_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout458_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout459_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout460_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout461_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout462_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout463_A (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout464_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout466_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout467_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout468_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout469_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout470_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout471_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout472_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout474_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout475_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout476_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout477_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout478_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout479_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout480_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout481_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout483_A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout484_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout485_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout486_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout487_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout488_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout489_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout490_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout491_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout492_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout493_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout494_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout495_A (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout496_A (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout497_A (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout498_A (.DIODE(net499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout500_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout501_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout502_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout503_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout504_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout505_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout506_A (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout507_A (.DIODE(net508));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout509_A (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout510_A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout511_A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout512_A (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout513_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout514_A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout515_A (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout516_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout523_A (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout526_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout527_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout528_A (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout531_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout532_A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout533_A (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout534_A (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout535_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout536_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout537_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout538_A (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout86_A (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout87_A (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout88_A (.DIODE(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout89_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout90_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout92_A (.DIODE(\u_usb_host.u_core._097_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout93_A (.DIODE(\u_usb_host.u_core._097_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout95_A (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout97_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0475_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout98_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0458_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout99_A (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold121_A (.DIODE(\u_usb_host.u_core.u_sie.data_ready_w ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold122_A (.DIODE(\u_usb_host.u_core.u_sie.data_idx_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold22_A (.DIODE(\u_usb_host.u_core.u_sie.data_idx_i ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold2_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(reg_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(reg_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(reg_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(reg_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(reg_cs));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(reg_wdata[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(reg_wdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(reg_wdata[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(reg_wdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(reg_wdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(cfg_cska_usb[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(reg_wdata[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(reg_wdata[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(reg_wdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(reg_wdata[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(reg_wdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(reg_wdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(reg_wdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(reg_wdata[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(reg_wdata[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(reg_wdata[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(cfg_cska_usb[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(reg_wdata[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(reg_wdata[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(reg_wdata[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(reg_wdata[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(reg_wdata[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(reg_wdata[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(reg_wdata[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(reg_wdata[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(reg_wdata[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(reg_wdata[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(cfg_cska_usb[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(reg_wdata[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(reg_wdata[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(reg_wdata[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(reg_wr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(usb_in_dn));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(usb_in_dp));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(usb_rstn));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(wbd_clk_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(cfg_cska_usb[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(reg_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(reg_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(reg_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(reg_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(reg_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_output48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_output60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_output74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_output75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._14__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._19__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._20__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._21__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._22__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._31__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._32__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._33__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._34__A_N  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._35__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._36__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._39__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._40__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._41__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._42__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._47__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._48__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._49__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._50__A_N  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._51__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._52__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._53__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._54__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._55__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._56__A_N  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb._57__A  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._043__A  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._044__A  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._048__A  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._048__B  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._049__A  (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._049__B  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._068__A  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._069__A  (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._070__A  (.DIODE(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._088__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._088__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._089__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._089__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._090__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._090__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._091__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._091__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._092__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._092__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._093__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._093__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._094__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._094__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._095__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._095__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._096__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._096__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._097__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._097__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._098__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._098__S1  (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._099__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._099__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._100__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._100__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._101__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._101__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._102__S0  (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._102__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._103__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._103__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._104__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._104__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._105__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._105__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._106__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._106__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._107__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._107__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._108__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._108__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._109__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._109__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._110__S0  (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._110__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._111__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._111__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._116__S0  (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._116__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._117__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._117__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._118__S0  (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._118__S1  (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._119__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._119__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._120__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._120__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._121__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._121__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._122__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._122__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._123__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._123__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._124__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._124__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._125__S0  (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._125__S1  (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._126__S0  (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._126__S1  (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._140__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._141__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._141__D  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._143__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._143__D  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._144__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._145__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._147__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._148__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._151__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._151__D  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._152__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._152__D  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._153__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._155__D  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._157__D  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._163__D  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._182__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._183__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._184__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._184__D  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._186__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._186__D  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._187__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._188__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._190__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._191__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._194__D  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._195__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._195__D  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._196__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._198__D  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._200__D  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._206__D  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._227__D  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._229__D  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._237__D  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._238__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._238__D  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._241__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._241__D  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._242__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._243__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._243__D  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._249__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._249__D  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._250__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._251__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._252__CLK  (.DIODE(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._260__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._261__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._262__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._272__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._273__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._273__D  (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._275__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._275__D  (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._276__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._277__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._279__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._280__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._283__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._283__D  (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._284__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._284__D  (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._285__CLK  (.DIODE(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._287__D  (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._289__D  (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._295__D  (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._312__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._313__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_cmd_if._314__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._021__A  (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._025__B  (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._033__A  (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._035__A1  (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._038__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._039__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._040__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._041__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._042__S  (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._043__S  (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._044__S  (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._045__S  (.DIODE(net569));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._046__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._047__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._048__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._049__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._051__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._052__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._053__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._056__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._058__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._062__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._063__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._064__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._065__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._066__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._067__S  (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._069__S  (.DIODE(net526));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._074__B  (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._151__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._152__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._161__GATE  (.DIODE(\u_usb_host.u_async_wb.u_resp_if._000_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_async_wb.u_resp_if._162__GATE  (.DIODE(\u_usb_host.u_async_wb.u_resp_if._001_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._209__A  (.DIODE(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._218__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._221__B  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._228__B  (.DIODE(\u_usb_host.u_core._003_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._243__A2  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._243__B1  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._245__A2  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._248__A  (.DIODE(\u_usb_host.reg_addr[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._249__B  (.DIODE(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._249__C_N  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._251__A  (.DIODE(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._252__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._252__B  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._255__C  (.DIODE(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._255__D  (.DIODE(\u_usb_host.reg_addr[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._257__A  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._258__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._258__B  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._259__B  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._260__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._260__B  (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._261__B  (.DIODE(\u_usb_host.reg_addr[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._263__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._263__B  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._264__B  (.DIODE(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._265__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._265__B  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._267__B  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._268__B  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._269__B  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._270__B  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._279__A  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._281__A  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._304__A  (.DIODE(\u_usb_host.u_core.usb_xfer_token_in_out_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._305__A  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ack_out_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._306__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._307__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._308__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._309__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._311__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._312__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._313__B  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._322__A0  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._323__A0  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._324__A0  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._326__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ack_out_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._326__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._326__B1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._327__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._328__B1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._329__A1  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._329__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._330__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._330__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._330__B1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._332__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._332__B1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._334__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._335__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._337__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._340__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._342__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._344__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__B1  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._346__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._347__A2  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._347__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._349__A2  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._349__B1  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._351__A2  (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._351__B1  (.DIODE(\u_usb_host.u_core._130_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._352__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._352__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._353__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._353__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._353__B1  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._353__B2  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._354__A2  (.DIODE(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._355__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._355__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._356__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._356__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._356__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._357__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._357__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._358__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._358__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._359__A2  (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._359__B1  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._359__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._360__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._361__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._361__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._362__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._362__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._362__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._363__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._363__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._364__A2  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._364__B1  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._365__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._365__B1  (.DIODE(\u_usb_host.u_core._130_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._366__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._366__B1  (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._367__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._367__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._368__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._368__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._369__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._369__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._369__B1  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._370__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._370__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._371__A2  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._371__B1  (.DIODE(\u_usb_host.u_core._130_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._372__A2  (.DIODE(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._372__B1  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._373__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.data_o[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._373__A2  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._373__B1  (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._374__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._375__A1  (.DIODE(\u_usb_host.u_core.usb_xfer_token_in_out_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._375__A2  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._375__B1  (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._376__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._377__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._378__A2  (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._379__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._381__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._383__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._385__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._386__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._387__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._388__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._389__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._390__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._391__B1  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._392__A2  (.DIODE(net87));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._395__B  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._397__A  (.DIODE(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._397__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._398__A  (.DIODE(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._398__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._399__A  (.DIODE(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._399__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._400__A  (.DIODE(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._400__B  (.DIODE(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._401__A  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._401__C  (.DIODE(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._402__A  (.DIODE(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._402__B  (.DIODE(\u_usb_host.u_core._033_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._427__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._428__D  (.DIODE(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._429__D  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._430__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._431__D  (.DIODE(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._432__D  (.DIODE(\u_usb_host.reg_wdata[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._433__D  (.DIODE(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._434__D  (.DIODE(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._436__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._436__D  (.DIODE(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._436__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._437__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._437__D  (.DIODE(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._438__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._438__D  (.DIODE(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._439__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._439__D  (.DIODE(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._440__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._440__D  (.DIODE(\u_usb_host.reg_wdata[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._441__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._441__D  (.DIODE(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._442__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._442__D  (.DIODE(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._443__CLK  (.DIODE(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._443__D  (.DIODE(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._444__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._445__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._446__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._447__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._448__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._449__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._450__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._451__CLK  (.DIODE(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._452__D  (.DIODE(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._489__D  (.DIODE(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._489__RESET_B  (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._490__D  (.DIODE(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._492__D  (.DIODE(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._500__RESET_B  (.DIODE(net372));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._508__D  (.DIODE(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._509__D  (.DIODE(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._510__D  (.DIODE(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._511__D  (.DIODE(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._512__D  (.DIODE(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._514__D  (.DIODE(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._515__D  (.DIODE(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._516__D  (.DIODE(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._517__D  (.DIODE(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._518__D  (.DIODE(\u_usb_host.reg_wdata[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._519__D  (.DIODE(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._520__D  (.DIODE(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._521__D  (.DIODE(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._522__D  (.DIODE(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._524__RESET_B  (.DIODE(net416));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._536__D  (.DIODE(\u_usb_host.u_core._003_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._550__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._551__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._552__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._556__D  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._564__D  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._567__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._568__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._569__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._576__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._577__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._578__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._579__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._580__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._581__GATE  (.DIODE(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._582__GATE  (.DIODE(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._583__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._585__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._586__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._587__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._588__GATE  (.DIODE(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._595__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._596__GATE  (.DIODE(\u_usb_host.u_core._033_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core._598__GATE  (.DIODE(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0796__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0797__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0799__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0803__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0804__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0804__B  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0806__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0807__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0807__B  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0811__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0811__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0813__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0813__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0815__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0815__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0817__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0817__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0819__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0821__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0821__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0822__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0822__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0824__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0824__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0826__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0826__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0828__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0828__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0830__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0830__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0831__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0832__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0834__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0834__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0836__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0837__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0838__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0838__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0839__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0839__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0840__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0840__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0841__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0841__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0843__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0843__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0844__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0844__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0844__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0845__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0845__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0846__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0846__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0847__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0847__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0848__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0848__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0849__A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0849__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0850__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0851__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0852__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0852__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0853__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0853__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0854__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0855__A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0855__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0856__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0458_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0856__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0857__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0458_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0857__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0858__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0858__B  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0860__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx.pop_i ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0861__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0861__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0862__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0862__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0863__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0863__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0863__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0864__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0864__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0865__A  (.DIODE(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0865__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0867__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0867__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0868__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0868__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0869__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0869__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0870__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0870__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0871__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0872__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0872__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0873__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0873__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0874__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0874__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0874__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0875__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0875__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0876__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0876__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0877__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0877__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0878__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0878__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0879__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0879__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0880__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0880__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0881__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0881__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0882__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0882__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0883__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0883__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0884__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0884__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0885__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0885__B  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0886__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0886__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0475_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0887__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0887__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0888__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0888__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0889__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0889__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0890__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0890__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0891__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0891__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0892__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0892__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0893__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0893__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0894__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0894__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0895__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0895__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0896__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0896__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0898__A0  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0898__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0903__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0903__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0909__A1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0909__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0912__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0913__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0917__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0918__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0920__A3  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0920__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0921__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0924__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0927__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0930__A1  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0930__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0932__A2  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0932__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0933__A2  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0936__A  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0936__B  (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0937__A2  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0938__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0939__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0940__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0942__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0944__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0944__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0945__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0946__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0948__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0951__A  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0951__B  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0952__A  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0952__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0954__A  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0954__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0957__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0957__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0959__A  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0961__B  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0963__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0965__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0966__A  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0966__B  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0967__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0968__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0969__A  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0969__B  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0970__A  (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0970__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0525_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0971__A  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0971__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0974__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0975__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0976__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0976__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0978__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0978__B  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0979__A  (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0979__B  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0980__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0980__C  (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0981__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0983__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0985__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0986__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0986__B  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0987__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0988__B  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0989__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0989__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0990__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0991__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0992__A  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0992__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0527_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0993__B  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0994__A  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0995__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._0998__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1001__A  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1001__B  (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1002__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1003__B  (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1005__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1005__B  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1007__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1009__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1009__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0575_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1010__A  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1010__B  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1011__A  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1011__B  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1012__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1014__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1014__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1016__C  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1017__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1018__A  (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1018__B  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1019__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1022__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1023__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1024__A  (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1024__B  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1025__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1026__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1027__A3  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1033__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1034__A3  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1039__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1045__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0610_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1045__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0611_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1050__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1052__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0618_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1054__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1055__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1056__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1057__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1058__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1059__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1060__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1060__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1064__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1065__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1065__C  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1066__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1067__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1068__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1069__B  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1070__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1071__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1072__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1073__C  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1074__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1076__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1077__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1078__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1078__C  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1079__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1080__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1083__B  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1083__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1084__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1085__C  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1089__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1090__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1091__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1091__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1092__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1099__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1100__A3  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1105__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1111__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0676_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1116__A2  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1116__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1119__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0684_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1120__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1121__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1123__B  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1123__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1124__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1127__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1128__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1129__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1129__C  (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1130__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1131__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1133__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1134__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1135__B  (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1136__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1137__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1139__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1140__C  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1141__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1143__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1145__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1148__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1151__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1152__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1155__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1156__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1157__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1158__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1159__A3  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1165__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1166__A3  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1171__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1182__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1184__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0102_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1184__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0113_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1185__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0114_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1186__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1187__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1189__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1190__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1193__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1193__C  (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1194__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1195__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1195__C  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1196__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1197__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1199__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1200__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1201__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1202__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1203__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1203__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1204__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1205__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1207__B  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1207__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1209__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1211__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1212__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1215__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1218__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1219__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1220__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1223__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1224__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1225__A3  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1231__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1232__A3  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1237__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1243__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0170_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1243__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0171_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1248__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1250__A  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0167_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1250__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1251__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0179_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1253__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1253__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1254__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1255__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1258__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1261__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1261__C  (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1262__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1263__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1264__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1266__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1267__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1269__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1270__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1271__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1272__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1273__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1274__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1275__B  (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1278__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1282__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1284__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1285__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1287__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1288__C  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1289__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1290__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1291__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1292__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1298__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1299__A3  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1304__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1315__A2  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1315__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1317__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0238_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1318__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0245_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1319__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1319__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1320__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1321__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1323__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1324__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1328__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1330__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1331__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1333__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1334__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1335__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1336__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1337__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1337__C  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1338__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1339__B  (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1339__C  (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1343__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1344__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1349__B  (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1352__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1354__C  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1356__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1357__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1358__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1359__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1365__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1366__A3  (.DIODE(net279));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1371__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1382__A2  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1382__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1384__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0304_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1385__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0311_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1386__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1387__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1388__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1389__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1390__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1391__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1395__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1397__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1400__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1401__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1402__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1403__C  (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1404__B  (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1404__C  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1405__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1406__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1410__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1411__B  (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1416__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0504_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1419__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1420__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1421__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1422__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1423__B  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1423__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1424__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0571_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1425__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1426__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1432__A2  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1432__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1433__A2  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1433__A3  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1438__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1449__A2  (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1449__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1451__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0370_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1452__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0377_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1453__B  (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1453__C  (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1454__C  (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1455__C  (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1457__C  (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1458__B  (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1462__C  (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1464__C  (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1465__C  (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1467__C  (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1468__C  (.DIODE(net296));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1469__B  (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1470__C  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0531_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1471__C  (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1472__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1473__C  (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1474__C  (.DIODE(net282));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1476__C  (.DIODE(net276));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1477__B  (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1478__B  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1478__C  (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1481__B  (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1484__C  (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1485__C  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1486__C  (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1487__B  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0504_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1490__C  (.DIODE(net280));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1491__B1  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1498__A2  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1498__A3  (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1499__A2  (.DIODE(net357));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1499__A3  (.DIODE(net278));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1504__A2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1515__A3  (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1517__D  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0441_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1518__B2  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0442_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1519__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1520__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1521__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1522__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1523__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1524__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1525__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1526__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1527__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1529__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1530__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1531__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1532__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1533__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1534__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1535__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1536__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1537__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1538__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1539__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1540__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1541__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1542__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1543__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1544__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1545__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1546__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1547__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1549__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1550__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1551__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1553__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1554__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1555__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1556__D  (.DIODE(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1557__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1558__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1559__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1560__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1561__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1562__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1563__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1565__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1566__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1567__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1568__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1569__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1570__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1571__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1572__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1573__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1574__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1575__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1576__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1577__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1578__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1579__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1580__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1581__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1582__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1583__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1584__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1585__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1586__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1587__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1588__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1589__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1590__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1591__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1593__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1594__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1595__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1596__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1597__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1598__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1599__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1600__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1601__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1602__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1603__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1604__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1605__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1606__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1607__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1609__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1610__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1611__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1612__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1613__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1614__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1615__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1616__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1617__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1618__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1619__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1620__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1621__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1622__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1623__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1624__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1625__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1626__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1627__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1628__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1629__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1630__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1631__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1632__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1633__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1634__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1635__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1636__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1637__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1638__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1639__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1640__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1641__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1642__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1643__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1644__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1645__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1646__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1647__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1648__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1649__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1650__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1651__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1652__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1653__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1654__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1655__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1656__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1657__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1658__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1659__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1660__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1661__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1662__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1663__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1664__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1665__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1666__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1667__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1668__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1669__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1670__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1671__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1672__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1673__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1674__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1675__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1676__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1677__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1678__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1679__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1680__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1681__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1682__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1683__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1684__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1685__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1686__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1687__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1688__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1689__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1690__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1691__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1692__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1693__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1694__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1695__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1696__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1697__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1698__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1699__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1700__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1701__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1702__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1703__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1704__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1705__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1706__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1707__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1708__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1709__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1710__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1711__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1712__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1713__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1714__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1715__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1717__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1718__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1719__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1720__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1721__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1722__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1723__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1724__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1725__D  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1726__D  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1727__D  (.DIODE(net175));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1728__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1729__D  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1730__D  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1731__D  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1732__D  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1733__D  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1734__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1735__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1736__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1737__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1738__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1739__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1740__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1741__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1742__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1743__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1744__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1745__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1746__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1747__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1748__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1749__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1750__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1751__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1752__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1753__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1754__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1755__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1757__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1758__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1759__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1760__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1761__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1762__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1763__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1764__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1765__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1766__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1767__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1768__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1769__D  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1770__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1771__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1773__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1774__D  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1775__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1776__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1777__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1778__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1779__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1780__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1781__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1782__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1783__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1784__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1785__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1786__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1787__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1788__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1789__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1790__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1791__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1792__D  (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1793__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1794__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1795__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1796__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1797__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1798__D  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1799__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1800__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1801__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1802__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1803__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1804__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1805__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1806__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1807__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1808__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1809__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1810__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1811__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1812__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1813__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1814__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1815__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1816__D  (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1817__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1818__D  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1819__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1820__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1821__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1822__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1823__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1824__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1825__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1826__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1827__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1828__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1829__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1830__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1831__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1832__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1833__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1834__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1835__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1836__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1837__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1838__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1839__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1840__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1841__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1842__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1843__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1844__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1845__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1846__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1847__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1848__D  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1849__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1850__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1851__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1852__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1853__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1854__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1862__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1863__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1864__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1865__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1866__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1867__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1868__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1869__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1871__RESET_B  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1876__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1877__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1878__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1879__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1880__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1881__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1882__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1883__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1884__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1885__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1886__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1887__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1888__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1889__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1890__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1891__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1892__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1893__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1894__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1895__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1896__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1897__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1898__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1899__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1900__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1901__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1902__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1903__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1904__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1905__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1906__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1907__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1931__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1933__CLK  (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1933__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0044_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1957__CLK  (.DIODE(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1964__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_rx._0075_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1975__D  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1976__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1977__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1978__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1979__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1980__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1981__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1982__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1983__D  (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1984__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1985__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1986__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1987__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1988__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1989__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1990__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1991__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1993__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1994__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1995__D  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1996__D  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1997__D  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1998__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._1999__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2000__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2001__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2002__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2003__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2004__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2005__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2006__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2007__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2008__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2009__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2010__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2011__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2012__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2013__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2014__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2015__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2016__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2017__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2018__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2019__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2020__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2021__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2022__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2023__D  (.DIODE(net180));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2024__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2025__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2026__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2027__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2028__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2029__D  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2030__D  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2031__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2032__D  (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2033__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2034__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2035__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2036__D  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2037__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2038__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2039__D  (.DIODE(net176));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2040__D  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2041__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2042__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2043__D  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2044__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2045__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2046__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2047__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2048__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2049__D  (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2050__D  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2051__D  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2052__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2053__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2054__D  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2055__D  (.DIODE(net177));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2056__D  (.DIODE(net167));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2057__D  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2058__D  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2059__D  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2060__D  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2061__D  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2062__D  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2063__D  (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2064__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2065__D  (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2066__D  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2067__D  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2068__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2069__D  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2070__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2071__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2072__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2073__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2074__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2075__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2076__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2077__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2078__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2079__D  (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2080__D  (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2081__D  (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2082__D  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2083__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2084__D  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2085__D  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2086__D  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2087__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2088__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2089__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2090__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2091__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2092__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2093__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2094__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2095__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2096__D  (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2097__D  (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2098__D  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2099__D  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2100__D  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2101__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2102__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2103__D  (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2104__D  (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2105__D  (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2106__D  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2107__D  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2108__D  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2109__D  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_rx._2110__D  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0796__A  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0796__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0797__A  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0797__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0799__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0799__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0803__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0804__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0804__B  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0806__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0807__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0807__B  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0811__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0811__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0813__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0813__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0815__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0815__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0819__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0819__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0821__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0821__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0822__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0822__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0824__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0824__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0826__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0826__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0828__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0828__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0832__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0834__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0834__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0836__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0836__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0837__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0837__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0838__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0838__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0839__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0839__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0840__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0841__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0841__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0843__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0844__C  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0845__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0846__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0846__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0847__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0847__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0475_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0848__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0848__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0849__A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0849__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0850__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0850__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0851__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0851__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0852__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0852__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0853__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0853__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0854__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0855__A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0856__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0857__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0858__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0858__B  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0860__B1  (.DIODE(\u_usb_host.u_core.fifo_tx_pop_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0861__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0862__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0865__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0867__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0868__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0869__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0870__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0873__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0462_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0873__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0874__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0463_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0875__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0454_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0875__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0876__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0876__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0877__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0473_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0877__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0878__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0452_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0878__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0879__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0465_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0879__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0880__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0880__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0881__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0881__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0882__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0882__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0883__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0884__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0884__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0885__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0885__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0886__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0886__B  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0887__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0472_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0887__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0889__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0466_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0889__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0890__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0467_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0890__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0891__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0892__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0468_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0892__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0893__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0457_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0893__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0894__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0895__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0469_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0895__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0930__A1  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0939__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0940__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0942__C  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0944__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0944__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0945__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0946__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0449_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0948__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0951__A  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0951__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0952__A  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0952__B  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0954__A  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0954__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0957__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0959__A  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0959__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0525_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0961__A  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0961__B  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0963__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0965__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0966__A  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0966__B  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0967__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0968__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0968__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0969__A  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0969__B  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0970__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0525_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0971__A  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0971__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0974__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0975__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0976__A  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0976__B  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0978__A  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0978__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0544_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0979__A  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0979__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0544_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0980__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0980__C  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0981__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0983__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0984__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0985__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0986__A  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0986__B  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0987__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0988__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0989__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0990__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0992__A  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0992__B  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0993__B  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0994__A  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0994__B  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0997__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._0998__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1000__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1000__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1001__A  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1001__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1002__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1003__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1005__A  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1005__B  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1009__A  (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1009__B  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1010__A  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1010__B  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1011__A  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1011__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1012__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1014__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1015__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1016__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1017__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1018__A  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1018__B  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1019__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1020__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1023__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1024__B  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1025__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1034__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1038__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1040__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0603_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1050__A2  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1050__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1052__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0612_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1052__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0618_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1055__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1056__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1057__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1059__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1060__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1063__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1064__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1065__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1065__C  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1066__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1067__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1068__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1068__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1069__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1070__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1073__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1074__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1076__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1078__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1080__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1080__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1081__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1082__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1083__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1085__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1086__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1086__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1089__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1090__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1091__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1093__A3  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1100__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1104__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1106__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0668_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1118__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0677_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1118__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0683_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1121__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1122__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1124__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1124__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1127__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1128__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1129__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1129__C  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1130__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1134__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1135__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1136__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1137__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1140__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1141__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1142__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1142__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1143__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1144__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1145__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1146__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1146__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1147__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1148__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1149__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1150__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1151__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1152__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1156__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1157__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1165__A3  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1166__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1170__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1172__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0098_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1182__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1184__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0113_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1186__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1187__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1188__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1190__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1190__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1193__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1194__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1195__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1195__C  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1196__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1199__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1200__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1201__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1202__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1206__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1207__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1208__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1208__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1209__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1210__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1213__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1214__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1215__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1216__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1217__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1218__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1219__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1220__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1223__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1232__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1236__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1238__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0163_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1248__A2  (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1248__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1250__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0172_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1250__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0178_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1252__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1254__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1254__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1255__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1256__B  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1258__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1261__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1261__C  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1262__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1264__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1265__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1266__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1267__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1267__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1269__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1270__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1271__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1273__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1275__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1277__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1278__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1280__B  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1281__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1283__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1283__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1284__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1285__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1286__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1288__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1290__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1291__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1298__A3  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1299__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1300__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0227_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1303__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1305__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0229_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1315__A2  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1315__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1317__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0238_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1320__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1320__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1321__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1322__B  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1324__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1328__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1329__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1331__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1332__B  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1333__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1334__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1334__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1335__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1336__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1337__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0516_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1337__C  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1338__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1339__B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1340__B  (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1342__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1344__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1346__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1347__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1347__C  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1349__B  (.DIODE(net274));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1350__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1351__B  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1351__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1352__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1354__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1357__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1358__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1365__A3  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1366__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1370__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1382__A2  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1382__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1383__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0287_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1384__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0304_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1387__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1387__C  (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1388__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1389__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1391__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1395__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1396__C  (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1398__B  (.DIODE(net240));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1399__B  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1400__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1401__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1401__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1402__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1403__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1404__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0516_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1404__C  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1405__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1406__B  (.DIODE(net273));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1409__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1411__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1413__B  (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1413__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1414__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1414__C  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1416__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0504_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1417__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1418__B  (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1418__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1419__C  (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1421__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1424__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1425__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1432__A3  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1433__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1437__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1449__A2  (.DIODE(net237));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1449__A3  (.DIODE(net197));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1450__A  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0353_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1451__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0370_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1454__B  (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1455__C  (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1456__B  (.DIODE(net239));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1458__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1458__C  (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1462__C  (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1463__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1467__C  (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1468__B  (.DIODE(net244));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1468__C  (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1469__B  (.DIODE(net232));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1470__C  (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1471__B  (.DIODE(net243));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1471__C  (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1473__C  (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1474__C  (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1475__C  (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1477__B  (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1479__C  (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1480__B  (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1482__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1482__C  (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1483__B  (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1483__C  (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1484__C  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0575_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1485__C  (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1487__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0504_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1488__B  (.DIODE(net250));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1489__C  (.DIODE(net198));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1490__C  (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1492__A3  (.DIODE(net194));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1499__A3  (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1503__A2  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1515__A2  (.DIODE(net238));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1517__B  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0435_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1517__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0441_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1519__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1520__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1521__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1522__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1523__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1524__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1525__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1526__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1527__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1528__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1529__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1530__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1531__D  (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1533__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1534__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1535__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1536__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1537__D  (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1538__D  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1539__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1540__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1541__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1542__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1543__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1544__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1545__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1546__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1547__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1549__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1550__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1551__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1552__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1553__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1554__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1555__D  (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1557__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1558__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1559__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1560__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1561__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1562__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1563__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1565__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1566__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1567__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1568__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1569__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1570__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1571__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1572__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1573__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1574__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1575__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1576__D  (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1577__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1578__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1579__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1581__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1582__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1583__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1584__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1585__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1586__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1587__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1588__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1589__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1590__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1591__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1592__D  (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1593__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1594__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1595__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1597__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1598__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1599__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1600__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1601__D  (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1602__D  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1603__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1604__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1605__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1606__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1607__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1608__D  (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1609__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1610__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1611__D  (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1613__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1614__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1615__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1616__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1617__D  (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1618__D  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1619__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1620__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1621__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1622__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1623__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1624__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1625__D  (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1626__D  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1627__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1628__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1629__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1630__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1631__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1632__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1633__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1634__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1635__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1637__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1638__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1639__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1640__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1641__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1642__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1643__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1644__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1645__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1646__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1647__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1648__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1649__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1650__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1651__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1652__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1653__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1654__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1655__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1656__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1657__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1658__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1659__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1660__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1661__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1662__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1663__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1664__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1665__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1666__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1667__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1668__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1669__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1670__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1671__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1672__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1673__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1674__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1675__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1676__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1677__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1678__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1679__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1680__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1681__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1682__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1683__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1684__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1685__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1686__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1687__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1688__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1689__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1690__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1691__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1692__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1693__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1694__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1695__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1696__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1697__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1698__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1699__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1701__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1702__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1703__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1704__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1705__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1706__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1707__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1708__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1709__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1710__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1711__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1712__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1713__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1714__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1715__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1716__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1717__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1718__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1719__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1720__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1721__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1722__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1723__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1724__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1725__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1726__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1727__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1728__D  (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1729__D  (.DIODE(net501));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1730__D  (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1731__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1732__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1733__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1734__D  (.DIODE(net458));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1735__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1736__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1737__D  (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1738__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1739__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1740__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1741__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1742__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1743__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1744__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1745__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1746__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1747__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1748__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1749__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1750__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1751__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1752__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1753__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1754__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1755__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1756__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1757__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1758__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1759__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1760__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1761__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1762__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1763__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1764__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1765__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1766__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1767__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1768__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1769__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1770__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1771__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1773__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1774__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1775__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1776__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1777__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1778__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1779__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1780__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1781__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1782__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1783__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1784__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1785__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1786__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1787__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1788__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1789__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1790__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1791__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1792__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1793__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1794__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1795__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1797__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1798__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1799__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1800__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1801__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1802__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1803__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1804__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1805__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1806__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1807__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1808__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1809__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1810__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1811__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1812__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1813__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1814__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1815__D  (.DIODE(net520));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1816__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1817__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1818__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1819__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1821__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1822__D  (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1823__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1824__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1825__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1826__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1827__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1828__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1829__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1830__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1831__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1832__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1833__D  (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1834__D  (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1835__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1836__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1837__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1838__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1839__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1840__D  (.DIODE(net513));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1841__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1842__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1843__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1844__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1845__D  (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1846__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1847__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1848__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1849__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1850__D  (.DIODE(net498));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1851__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1852__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1853__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1854__D  (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1857__RESET_B  (.DIODE(net367));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1862__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1863__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1864__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1865__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1866__D  (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1867__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1868__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1869__D  (.DIODE(net464));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1870__RESET_B  (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1871__RESET_B  (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1872__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1873__RESET_B  (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1874__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1875__RESET_B  (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1876__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1877__D  (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1878__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1879__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1880__D  (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1881__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1882__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1883__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1884__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1885__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1886__D  (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1887__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1888__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1889__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1890__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1891__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1892__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1893__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1894__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1895__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1896__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1897__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1898__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1899__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1900__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1901__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1902__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1903__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1904__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1905__D  (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1906__D  (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1907__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1908__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0019_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1923__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0034_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1932__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0043_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1933__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0044_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1941__CLK  (.DIODE(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1950__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0061_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1952__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0063_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1963__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0074_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1964__GATE  (.DIODE(\u_usb_host.u_core.u_fifo_tx._0075_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1969__CLK  (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1974__CLK  (.DIODE(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1975__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1976__D  (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1977__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1978__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1979__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1980__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1981__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1982__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1983__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1984__D  (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1985__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1986__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1987__D  (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1988__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1989__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1990__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1991__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1992__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1993__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1994__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1995__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1997__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1998__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._1999__D  (.DIODE(net523));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2000__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2001__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2002__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2003__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2004__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2005__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2006__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2007__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2008__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2009__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2010__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2011__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2012__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2013__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2014__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2015__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2016__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2017__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2018__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2019__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2020__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2021__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2022__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2023__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2024__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2025__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2026__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2027__D  (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2028__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2029__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2030__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2031__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2032__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2033__D  (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2034__D  (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2035__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2036__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2037__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2038__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2039__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2040__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2041__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2042__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2043__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2044__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2045__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2046__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2047__D  (.DIODE(net517));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2048__D  (.DIODE(net510));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2049__D  (.DIODE(net500));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2050__D  (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2051__D  (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2052__D  (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2053__D  (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2054__D  (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2055__D  (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2056__D  (.DIODE(net511));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2057__D  (.DIODE(net503));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2058__D  (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2059__D  (.DIODE(net483));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2060__D  (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2061__D  (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2062__D  (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2063__D  (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2064__D  (.DIODE(net512));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2065__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2066__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2067__D  (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2068__D  (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2069__D  (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2070__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2071__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2072__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2073__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2074__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2075__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2076__D  (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2077__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2078__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2079__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2080__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2081__D  (.DIODE(net505));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2082__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2083__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2084__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2085__D  (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2086__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2087__D  (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2088__D  (.DIODE(net516));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2089__D  (.DIODE(net504));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2090__D  (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2091__D  (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2092__D  (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2093__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2094__D  (.DIODE(net461));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2095__D  (.DIODE(net522));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2096__D  (.DIODE(net514));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2097__D  (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2098__D  (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2099__D  (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2100__D  (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2101__D  (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2102__D  (.DIODE(net462));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2103__D  (.DIODE(\u_usb_host.u_core.u_fifo_tx.data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2104__D  (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2105__D  (.DIODE(net507));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2106__D  (.DIODE(net497));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2107__D  (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2108__D  (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2109__D  (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2110__D  (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2111__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2112__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2113__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2114__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2115__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_fifo_tx._2116__RESET_B  (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._331__B  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._344__B  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._350__A  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._351__B1  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._357__A  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._364__B  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._366__B  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._376__A  (.DIODE(\u_usb_host.u_core.u_sie.data_ready_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._378__B1  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._380__B  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._381__B  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._382__B  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._384__A2  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._391__A  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._409__A2  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._411__A  (.DIODE(\u_usb_host.u_core.u_sie.data_ready_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._412__B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._414__A  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._414__B  (.DIODE(\u_usb_host.u_core.u_sie._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._416__B  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._417__B1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._417__C1  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._421__A2  (.DIODE(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._421__B1  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._422__B  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._425__A1  (.DIODE(\u_usb_host.u_core.u_sie.data_ready_w ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._425__A2  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._426__B1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._427__A2  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._428__A2  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._432__B1  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._437__B  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._441__B  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._442__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._443__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._444__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._445__B  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._446__B  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._447__A1  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._464__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._465__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._466__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._467__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._468__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._469__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._470__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._471__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._498__A1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._498__B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._502__A1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._502__B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._506__A2  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._508__A2  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._508__B1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._512__A2  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._512__B1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._520__A1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._520__B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._524__A1  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._524__B1  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._528__A2  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._546__B1  (.DIODE(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._557__B  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._558__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._561__B  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._563__B  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._564__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._566__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._568__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._570__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._572__B1  (.DIODE(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._581__A1  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._581__A2  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._582__A2  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._582__B1  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._584__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._585__A1  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._586__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._586__A2  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._588__A2  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._589__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._589__C1  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._590__B  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._592__A2  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._592__B1  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._592__B2  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._593__S  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._595__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._596__A1  (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._596__B1  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._597__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._597__A2  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._599__A2  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._600__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._600__C1  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._601__B  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._603__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._603__A2  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._605__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._605__B1  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._608__A2  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._608__B1  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._608__B2  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._609__S  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._611__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._612__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._612__A2  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._614__A2  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._615__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._615__C1  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._616__B  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._619__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._619__A2  (.DIODE(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._620__B2  (.DIODE(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._621__S  (.DIODE(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._623__A2  (.DIODE(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._624__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._624__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._624__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._625__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._625__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._625__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._626__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._626__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._626__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._627__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._627__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._627__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._628__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._628__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._628__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._629__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._629__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._629__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._630__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._630__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._630__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._631__A0  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._631__A1  (.DIODE(\u_usb_host.u_core.fifo_tx_data_w[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._631__S  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._632__A  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._634__B  (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._635__C  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._650__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._651__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._652__RESET_B  (.DIODE(net403));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._675__RESET_B  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._678__RESET_B  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._696__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._697__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._700__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._701__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._702__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._703__RESET_B  (.DIODE(net384));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._704__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._705__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._706__D  (.DIODE(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._709__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._710__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._711__RESET_B  (.DIODE(net398));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._741__D  (.DIODE(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._755__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._756__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._757__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._758__D  (.DIODE(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._761__D  (.DIODE(\u_usb_host.u_core.u_sie._042_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._772__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._773__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._774__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._777__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._778__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._782__CLK  (.DIODE(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._783__GATE  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._791__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._792__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[1] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._793__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._794__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._795__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._796__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._797__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_core.u_sie._798__A  (.DIODE(\u_usb_host.u_core.u_sie.data_buffer_q[7] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._187__A  (.DIODE(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._195__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._211__A  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._212__B  (.DIODE(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._213__C  (.DIODE(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._214__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._221__C  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._229__C  (.DIODE(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._231__A  (.DIODE(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._232__A  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._234__C  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._235__A1  (.DIODE(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._237__A  (.DIODE(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._238__A  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._247__A1  (.DIODE(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._248__A1  (.DIODE(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._250__A  (.DIODE(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._255__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._266__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._266__B  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._268__B1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._269__A  (.DIODE(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._275__A1  (.DIODE(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._280__A1  (.DIODE(\u_usb_host.u_core.u_sie.utmi_data_o[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._280__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._282__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._284__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._286__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._288__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._290__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._292__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._295__B  (.DIODE(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._296__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._302__B1  (.DIODE(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._303__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._305__B1  (.DIODE(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._305__C1  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._318__B  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._333__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._336__B  (.DIODE(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._337__B  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._338__A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._343__A2  (.DIODE(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._345__B  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._349__A1  (.DIODE(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._350__A  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._351__A2  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._353__A2  (.DIODE(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._361__A1  (.DIODE(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._372__D  (.DIODE(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._372__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._387__SET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._388__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._389__RESET_B  (.DIODE(net409));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._391__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._392__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._393__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._394__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._395__RESET_B  (.DIODE(net395));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_phy._409__RESET_B  (.DIODE(net392));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._1__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst._2__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_usb_rst.u_buf.genblk1.u_mux_A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst._1__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst._2__RESET_B  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_usb_host.u_wb_rst.u_buf.genblk1.u_mux_A1  (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_A (.DIODE(usb_clk));
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_396 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_13 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_514 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_154 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_480 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_152 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_451 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_364 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_283 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_347 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_19 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_12 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_159 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_282 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_252 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_254 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_322 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_374 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_242 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_640 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_344 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_706 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_131 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_686 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_448 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_569 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_114 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_434 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_786 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_513 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_264 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_646 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_676 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_797 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_770 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_255 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_99 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_370 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_514 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_508 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_77 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_618 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_635 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_702 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_746 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_145 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_398 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_106 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_610 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_114 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_22 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_217 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_374 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_384 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_514 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_331 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_631 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_965 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_622 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_68 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_23 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_475 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_428 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_648 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_258 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_326 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_704 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_171 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_584 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_178 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_534 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_889 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_350 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_542 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_413 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_196 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_329 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_32 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_12 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_231 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_539 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_208 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_435 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_269 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_452 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_662 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_367 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_961 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_384 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_410 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_634 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_949 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_479 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_483 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_562 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_126 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_142 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_762 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_340 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_371 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_775 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_16 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_380 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_778 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_168 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_283 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_672 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_467 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_364 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_933 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_224 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_348 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_747 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_426 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_777 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_658 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_686 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_338 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_110 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_579 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_650 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_518 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_663 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_67 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_739 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_622 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_692 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_571 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_741 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_473 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_548 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_11 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_293 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_724 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_748 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_554 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_709 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_110 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_295 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_234 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_679 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_764 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1057 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_271 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_107 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_515 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_509 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_717 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_32 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_644 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_8 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_343 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_364 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1057 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_422 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_582 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_382 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_314 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_438 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_438 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_382 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_460 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_333 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_202 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_318 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_426 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_370 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_302 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_260 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_436 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_220 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_22 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_230 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_395 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_464 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_548 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_16 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_286 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_343 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_454 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_400 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_540 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_375 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_18 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_504 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1049 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_275 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_1 _01_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[0] ),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 _02_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[1] ),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_2 _03_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[2] ),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_2 _04_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[3] ),
    .X(net74));
 sky130_fd_sc_hd__clkbuf_2 _05_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[4] ),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 _06_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[5] ),
    .X(net76));
 sky130_fd_sc_hd__clkbuf_1 _07_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[6] ),
    .X(net77));
 sky130_fd_sc_hd__clkbuf_1 _08_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[7] ),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 _09_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[8] ),
    .X(net79));
 sky130_fd_sc_hd__and4bb_1 _0_ (.A_N(net11),
    .B_N(net13),
    .C(net14),
    .D(net12),
    .X(\u_usb_host.u_async_wb.wbm_cyc_i ));
 sky130_fd_sc_hd__clkbuf_1 _10_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[9] ),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 _11_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[10] ),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 _12_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[11] ),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_1 _13_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[12] ),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_1 _14_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[13] ),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 _15_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[14] ),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 _16_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[15] ),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_1 _17_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[16] ),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 _18_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[17] ),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 _19_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[18] ),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 _20_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[19] ),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 _21_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[20] ),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 _22_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[21] ),
    .X(net62));
 sky130_fd_sc_hd__clkbuf_1 _23_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[22] ),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 _24_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[23] ),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_1 _25_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[24] ),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_1 _26_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[25] ),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 _27_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[26] ),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 _28_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[27] ),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 _29_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[28] ),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_1 _30_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[29] ),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 _31_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[30] ),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 _32_ (.A(\u_usb_host.u_async_wb.u_resp_if.rd_data[31] ),
    .X(net73));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_app_clk (.A(app_clk),
    .X(clknet_0_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._171_  (.A(\u_usb_host.u_core._171_ ),
    .X(\clknet_0_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._172_  (.A(\u_usb_host.u_core._172_ ),
    .X(\clknet_0_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._178_  (.A(\u_usb_host.u_core._178_ ),
    .X(\clknet_0_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._183_  (.A(\u_usb_host.u_core._183_ ),
    .X(\clknet_0_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._184_  (.A(\u_usb_host.u_core._184_ ),
    .X(\clknet_0_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._185_  (.A(\u_usb_host.u_core._185_ ),
    .X(\clknet_0_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._186_  (.A(\u_usb_host.u_core._186_ ),
    .X(\clknet_0_u_usb_host.u_core._186_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._192_  (.A(\u_usb_host.u_core._192_ ),
    .X(\clknet_0_u_usb_host.u_core._192_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._193_  (.A(\u_usb_host.u_core._193_ ),
    .X(\clknet_0_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core._200_  (.A(\u_usb_host.u_core._200_ ),
    .X(\clknet_0_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0784_  (.A(\u_usb_host.u_core.u_fifo_rx._0784_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0785_  (.A(\u_usb_host.u_core.u_fifo_rx._0785_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0786_  (.A(\u_usb_host.u_core.u_fifo_rx._0786_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_rx._0787_  (.A(\u_usb_host.u_core.u_fifo_rx._0787_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_rx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0721_  (.A(\u_usb_host.u_core.u_fifo_tx._0721_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0722_  (.A(\u_usb_host.u_core.u_fifo_tx._0722_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0723_  (.A(\u_usb_host.u_core.u_fifo_tx._0723_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0724_  (.A(\u_usb_host.u_core.u_fifo_tx._0724_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0725_  (.A(\u_usb_host.u_core.u_fifo_tx._0725_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0726_  (.A(\u_usb_host.u_core.u_fifo_tx._0726_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0727_  (.A(\u_usb_host.u_core.u_fifo_tx._0727_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0728_  (.A(\u_usb_host.u_core.u_fifo_tx._0728_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0729_  (.A(\u_usb_host.u_core.u_fifo_tx._0729_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0730_  (.A(\u_usb_host.u_core.u_fifo_tx._0730_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0731_  (.A(\u_usb_host.u_core.u_fifo_tx._0731_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0732_  (.A(\u_usb_host.u_core.u_fifo_tx._0732_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0733_  (.A(\u_usb_host.u_core.u_fifo_tx._0733_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0734_  (.A(\u_usb_host.u_core.u_fifo_tx._0734_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0735_  (.A(\u_usb_host.u_core.u_fifo_tx._0735_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0736_  (.A(\u_usb_host.u_core.u_fifo_tx._0736_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0737_  (.A(\u_usb_host.u_core.u_fifo_tx._0737_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0738_  (.A(\u_usb_host.u_core.u_fifo_tx._0738_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0739_  (.A(\u_usb_host.u_core.u_fifo_tx._0739_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0740_  (.A(\u_usb_host.u_core.u_fifo_tx._0740_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0741_  (.A(\u_usb_host.u_core.u_fifo_tx._0741_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0742_  (.A(\u_usb_host.u_core.u_fifo_tx._0742_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0743_  (.A(\u_usb_host.u_core.u_fifo_tx._0743_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0744_  (.A(\u_usb_host.u_core.u_fifo_tx._0744_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0745_  (.A(\u_usb_host.u_core.u_fifo_tx._0745_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0746_  (.A(\u_usb_host.u_core.u_fifo_tx._0746_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0747_  (.A(\u_usb_host.u_core.u_fifo_tx._0747_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0748_  (.A(\u_usb_host.u_core.u_fifo_tx._0748_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0749_  (.A(\u_usb_host.u_core.u_fifo_tx._0749_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0750_  (.A(\u_usb_host.u_core.u_fifo_tx._0750_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0751_  (.A(\u_usb_host.u_core.u_fifo_tx._0751_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0752_  (.A(\u_usb_host.u_core.u_fifo_tx._0752_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0753_  (.A(\u_usb_host.u_core.u_fifo_tx._0753_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0754_  (.A(\u_usb_host.u_core.u_fifo_tx._0754_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0755_  (.A(\u_usb_host.u_core.u_fifo_tx._0755_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0756_  (.A(\u_usb_host.u_core.u_fifo_tx._0756_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0757_  (.A(\u_usb_host.u_core.u_fifo_tx._0757_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0758_  (.A(\u_usb_host.u_core.u_fifo_tx._0758_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0759_  (.A(\u_usb_host.u_core.u_fifo_tx._0759_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0760_  (.A(\u_usb_host.u_core.u_fifo_tx._0760_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0761_  (.A(\u_usb_host.u_core.u_fifo_tx._0761_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0762_  (.A(\u_usb_host.u_core.u_fifo_tx._0762_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0763_  (.A(\u_usb_host.u_core.u_fifo_tx._0763_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0764_  (.A(\u_usb_host.u_core.u_fifo_tx._0764_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0765_  (.A(\u_usb_host.u_core.u_fifo_tx._0765_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0766_  (.A(\u_usb_host.u_core.u_fifo_tx._0766_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0767_  (.A(\u_usb_host.u_core.u_fifo_tx._0767_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0768_  (.A(\u_usb_host.u_core.u_fifo_tx._0768_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0769_  (.A(\u_usb_host.u_core.u_fifo_tx._0769_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0770_  (.A(\u_usb_host.u_core.u_fifo_tx._0770_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0771_  (.A(\u_usb_host.u_core.u_fifo_tx._0771_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0772_  (.A(\u_usb_host.u_core.u_fifo_tx._0772_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0773_  (.A(\u_usb_host.u_core.u_fifo_tx._0773_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0774_  (.A(\u_usb_host.u_core.u_fifo_tx._0774_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0775_  (.A(\u_usb_host.u_core.u_fifo_tx._0775_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0776_  (.A(\u_usb_host.u_core.u_fifo_tx._0776_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0777_  (.A(\u_usb_host.u_core.u_fifo_tx._0777_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0778_  (.A(\u_usb_host.u_core.u_fifo_tx._0778_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0779_  (.A(\u_usb_host.u_core.u_fifo_tx._0779_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0780_  (.A(\u_usb_host.u_core.u_fifo_tx._0780_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0781_  (.A(\u_usb_host.u_core.u_fifo_tx._0781_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0782_  (.A(\u_usb_host.u_core.u_fifo_tx._0782_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0783_  (.A(\u_usb_host.u_core.u_fifo_tx._0783_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0784_  (.A(\u_usb_host.u_core.u_fifo_tx._0784_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0785_  (.A(\u_usb_host.u_core.u_fifo_tx._0785_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0786_  (.A(\u_usb_host.u_core.u_fifo_tx._0786_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_fifo_tx._0787_  (.A(\u_usb_host.u_core.u_fifo_tx._0787_ ),
    .X(\clknet_0_u_usb_host.u_core.u_fifo_tx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._294_  (.A(\u_usb_host.u_core.u_sie._294_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._294_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._295_  (.A(\u_usb_host.u_core.u_sie._295_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._295_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._296_  (.A(\u_usb_host.u_core.u_sie._296_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._296_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._305_  (.A(\u_usb_host.u_core.u_sie._305_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._305_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._306_  (.A(\u_usb_host.u_core.u_sie._306_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._307_  (.A(\u_usb_host.u_core.u_sie._307_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._307_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._308_  (.A(\u_usb_host.u_core.u_sie._308_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._308_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._310_  (.A(\u_usb_host.u_core.u_sie._310_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._310_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._311_  (.A(\u_usb_host.u_core.u_sie._311_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._311_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_core.u_sie._312_  (.A(\u_usb_host.u_core.u_sie._312_ ),
    .X(\clknet_0_u_usb_host.u_core.u_sie._312_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._173_  (.A(\u_usb_host.u_phy._173_ ),
    .X(\clknet_0_u_usb_host.u_phy._173_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._176_  (.A(\u_usb_host.u_phy._176_ ),
    .X(\clknet_0_u_usb_host.u_phy._176_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._178_  (.A(\u_usb_host.u_phy._178_ ),
    .X(\clknet_0_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._179_  (.A(\u_usb_host.u_phy._179_ ),
    .X(\clknet_0_u_usb_host.u_phy._179_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_0_u_usb_host.u_phy._182_  (.A(\u_usb_host.u_phy._182_ ),
    .X(\clknet_0_u_usb_host.u_phy._182_ ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_usb_clk (.A(net565),
    .X(clknet_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_app_clk (.A(clknet_0_app_clk),
    .X(clknet_1_0__leaf_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._171_  (.A(\clknet_0_u_usb_host.u_core._171_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._172_  (.A(\clknet_0_u_usb_host.u_core._172_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._178_  (.A(\clknet_0_u_usb_host.u_core._178_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._183_  (.A(\clknet_0_u_usb_host.u_core._183_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._184_  (.A(\clknet_0_u_usb_host.u_core._184_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._185_  (.A(\clknet_0_u_usb_host.u_core._185_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._186_  (.A(\clknet_0_u_usb_host.u_core._186_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._186_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._192_  (.A(\clknet_0_u_usb_host.u_core._192_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._192_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core._193_  (.A(\clknet_0_u_usb_host.u_core._193_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0784_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0785_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0786_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_rx._0787_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0784_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0785_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0786_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_fifo_tx._0787_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._294_  (.A(\clknet_0_u_usb_host.u_core.u_sie._294_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._294_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._295_  (.A(\clknet_0_u_usb_host.u_core.u_sie._295_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._296_  (.A(\clknet_0_u_usb_host.u_core.u_sie._296_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._305_  (.A(\clknet_0_u_usb_host.u_core.u_sie._305_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._307_  (.A(\clknet_0_u_usb_host.u_core.u_sie._307_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._307_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._308_  (.A(\clknet_0_u_usb_host.u_core.u_sie._308_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._308_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._310_  (.A(\clknet_0_u_usb_host.u_core.u_sie._310_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._311_  (.A(\clknet_0_u_usb_host.u_core.u_sie._311_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._311_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_core.u_sie._312_  (.A(\clknet_0_u_usb_host.u_core.u_sie._312_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._173_  (.A(\clknet_0_u_usb_host.u_phy._173_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._173_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._176_  (.A(\clknet_0_u_usb_host.u_phy._176_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._176_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._178_  (.A(\clknet_0_u_usb_host.u_phy._178_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._179_  (.A(\clknet_0_u_usb_host.u_phy._179_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._179_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_0__f_u_usb_host.u_phy._182_  (.A(\clknet_0_u_usb_host.u_phy._182_ ),
    .X(\clknet_1_0__leaf_u_usb_host.u_phy._182_ ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_app_clk (.A(clknet_0_app_clk),
    .X(clknet_1_1__leaf_app_clk));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._035_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._036_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._037_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_cmd_if._038_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._014_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._015_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._016_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_async_wb.u_resp_if._017_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._171_  (.A(\clknet_0_u_usb_host.u_core._171_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._172_  (.A(\clknet_0_u_usb_host.u_core._172_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._178_  (.A(\clknet_0_u_usb_host.u_core._178_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._183_  (.A(\clknet_0_u_usb_host.u_core._183_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._184_  (.A(\clknet_0_u_usb_host.u_core._184_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._185_  (.A(\clknet_0_u_usb_host.u_core._185_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._186_  (.A(\clknet_0_u_usb_host.u_core._186_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._186_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._192_  (.A(\clknet_0_u_usb_host.u_core._192_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._192_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core._193_  (.A(\clknet_0_u_usb_host.u_core._193_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0784_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0785_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0786_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_rx._0787_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0721_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0722_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0723_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0724_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0725_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0726_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0727_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0728_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0729_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0730_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0731_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0732_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0733_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0734_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0735_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0736_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0737_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0738_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0739_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0740_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0741_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0742_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0743_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0744_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0745_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0746_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0747_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0748_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0749_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0750_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0751_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0752_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0753_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0754_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0755_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0756_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0757_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0758_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0759_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0760_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0761_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0762_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0763_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0764_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0765_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0766_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0767_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0768_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0769_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0770_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0771_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0772_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0773_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0774_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0775_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0776_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0777_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0778_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0779_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0780_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0781_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0782_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0783_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0784_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0785_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0786_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_fifo_tx._0787_  (.A(\clknet_0_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._294_  (.A(\clknet_0_u_usb_host.u_core.u_sie._294_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._294_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._295_  (.A(\clknet_0_u_usb_host.u_core.u_sie._295_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._296_  (.A(\clknet_0_u_usb_host.u_core.u_sie._296_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._305_  (.A(\clknet_0_u_usb_host.u_core.u_sie._305_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._307_  (.A(\clknet_0_u_usb_host.u_core.u_sie._307_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._307_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._308_  (.A(\clknet_0_u_usb_host.u_core.u_sie._308_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._308_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._310_  (.A(\clknet_0_u_usb_host.u_core.u_sie._310_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._311_  (.A(\clknet_0_u_usb_host.u_core.u_sie._311_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._311_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_core.u_sie._312_  (.A(\clknet_0_u_usb_host.u_core.u_sie._312_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._173_  (.A(\clknet_0_u_usb_host.u_phy._173_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._173_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._176_  (.A(\clknet_0_u_usb_host.u_phy._176_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._176_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._178_  (.A(\clknet_0_u_usb_host.u_phy._178_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._179_  (.A(\clknet_0_u_usb_host.u_phy._179_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._179_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_1_1__f_u_usb_host.u_phy._182_  (.A(\clknet_0_u_usb_host.u_phy._182_ ),
    .X(\clknet_1_1__leaf_u_usb_host.u_phy._182_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_0__f_u_usb_host.u_core.u_sie._306_  (.A(\clknet_0_u_usb_host.u_core.u_sie._306_ ),
    .X(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_1__f_u_usb_host.u_core.u_sie._306_  (.A(\clknet_0_u_usb_host.u_core.u_sie._306_ ),
    .X(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_2__f_u_usb_host.u_core.u_sie._306_  (.A(\clknet_0_u_usb_host.u_core.u_sie._306_ ),
    .X(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._039_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._040_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._041_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_cmd_if._042_  (.A(\clknet_0_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_resp_if._018_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_async_wb.u_resp_if._019_  (.A(\clknet_0_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_core._200_  (.A(\clknet_0_u_usb_host.u_core._200_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__clkbuf_16 \clkbuf_2_3__f_u_usb_host.u_core.u_sie._306_  (.A(\clknet_0_u_usb_host.u_core.u_sie._306_ ),
    .X(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_0_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_0_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_1_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_1_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_2_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_2_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_3_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_3_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_4_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_4_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_5_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_5_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_6_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_6_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_3_7_0_usb_clk (.A(clknet_0_usb_clk),
    .X(clknet_3_7_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_usb_clk (.A(clknet_3_0_0_usb_clk),
    .X(clknet_leaf_0_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_10_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_11_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_12_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_13_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_14_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_15_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_16_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_17_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_18_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_18_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_19_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_usb_clk (.A(clknet_3_1_0_usb_clk),
    .X(clknet_leaf_1_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_20_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_21_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_22_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_23_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_24_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_25_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_26_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_27_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_27_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_28_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_29_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_usb_clk (.A(clknet_3_0_0_usb_clk),
    .X(clknet_leaf_2_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_30_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_usb_clk (.A(clknet_3_7_0_usb_clk),
    .X(clknet_leaf_31_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_32_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_34_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_35_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_36_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_37_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_usb_clk (.A(clknet_3_3_0_usb_clk),
    .X(clknet_leaf_38_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_39_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_3_usb_clk (.A(clknet_3_1_0_usb_clk),
    .X(clknet_leaf_3_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_usb_clk (.A(clknet_3_6_0_usb_clk),
    .X(clknet_leaf_40_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_42_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_43_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_44_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_usb_clk (.A(clknet_3_3_0_usb_clk),
    .X(clknet_leaf_45_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_usb_clk (.A(clknet_3_3_0_usb_clk),
    .X(clknet_leaf_46_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_usb_clk (.A(clknet_3_3_0_usb_clk),
    .X(clknet_leaf_47_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_49_usb_clk (.A(clknet_3_1_0_usb_clk),
    .X(clknet_leaf_49_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_usb_clk (.A(clknet_3_1_0_usb_clk),
    .X(clknet_leaf_4_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_usb_clk (.A(clknet_3_1_0_usb_clk),
    .X(clknet_leaf_51_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_53_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_54_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_55_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_56_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_57_usb_clk (.A(clknet_3_2_0_usb_clk),
    .X(clknet_leaf_57_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_usb_clk (.A(clknet_3_0_0_usb_clk),
    .X(clknet_leaf_58_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_59_usb_clk (.A(clknet_3_0_0_usb_clk),
    .X(clknet_leaf_59_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_5_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_6_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_7_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_usb_clk (.A(clknet_3_4_0_usb_clk),
    .X(clknet_leaf_8_usb_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_usb_clk (.A(clknet_3_5_0_usb_clk),
    .X(clknet_leaf_9_usb_clk));
 sky130_fd_sc_hd__buf_2 fanout100 (.A(net101),
    .X(net100));
 sky130_fd_sc_hd__buf_2 fanout101 (.A(\u_usb_host.u_core.u_sie._166_ ),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(\u_usb_host.u_core.u_fifo_tx._0475_ ),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_4 fanout103 (.A(\u_usb_host.u_core.u_fifo_tx._0458_ ),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_4 fanout104 (.A(\u_usb_host.u_core.u_fifo_tx._0456_ ),
    .X(net104));
 sky130_fd_sc_hd__buf_2 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_4 fanout106 (.A(\u_usb_host.u_core.u_sie._164_ ),
    .X(net106));
 sky130_fd_sc_hd__buf_2 fanout107 (.A(\u_usb_host.u_async_wb.s_cmd_rd_empty ),
    .X(net107));
 sky130_fd_sc_hd__clkbuf_2 fanout108 (.A(\u_usb_host.u_async_wb.s_cmd_rd_empty ),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_2 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_2 fanout110 (.A(\u_usb_host.u_async_wb.s_cmd_rd_empty ),
    .X(net110));
 sky130_fd_sc_hd__clkbuf_2 fanout111 (.A(\u_usb_host.u_core.u_sie._176_ ),
    .X(net111));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout112 (.A(\u_usb_host.u_core.u_sie._176_ ),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_2 fanout114 (.A(\u_usb_host.u_core.status_sie_idle_w ),
    .X(net114));
 sky130_fd_sc_hd__buf_2 fanout115 (.A(\u_usb_host.u_phy._065_ ),
    .X(net115));
 sky130_fd_sc_hd__buf_2 fanout116 (.A(\u_usb_host.u_phy._064_ ),
    .X(net116));
 sky130_fd_sc_hd__clkbuf_4 fanout117 (.A(\u_usb_host.u_phy._058_ ),
    .X(net117));
 sky130_fd_sc_hd__buf_2 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__clkbuf_2 fanout119 (.A(net126),
    .X(net119));
 sky130_fd_sc_hd__buf_2 fanout120 (.A(net121),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_2 fanout121 (.A(net126),
    .X(net121));
 sky130_fd_sc_hd__buf_2 fanout122 (.A(net126),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_2 fanout123 (.A(net126),
    .X(net123));
 sky130_fd_sc_hd__buf_2 fanout124 (.A(net125),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_2 fanout125 (.A(net126),
    .X(net125));
 sky130_fd_sc_hd__clkbuf_4 fanout126 (.A(\u_usb_host.u_core.fifo_rx_data_w[7] ),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_4 fanout127 (.A(net134),
    .X(net127));
 sky130_fd_sc_hd__buf_2 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net134),
    .X(net129));
 sky130_fd_sc_hd__buf_2 fanout130 (.A(net134),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 fanout131 (.A(net134),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net134),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_2 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__buf_4 fanout134 (.A(\u_usb_host.u_core.fifo_rx_data_w[6] ),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_4 fanout135 (.A(net137),
    .X(net135));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout136 (.A(net137),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_2 fanout137 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net138));
 sky130_fd_sc_hd__buf_2 fanout139 (.A(net142),
    .X(net139));
 sky130_fd_sc_hd__buf_2 fanout140 (.A(net142),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net142),
    .X(net141));
 sky130_fd_sc_hd__buf_2 fanout142 (.A(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_4 fanout143 (.A(net146),
    .X(net143));
 sky130_fd_sc_hd__buf_2 fanout144 (.A(net146),
    .X(net144));
 sky130_fd_sc_hd__buf_2 fanout145 (.A(net146),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_2 fanout146 (.A(\u_usb_host.u_core.fifo_rx_data_w[4] ),
    .X(net146));
 sky130_fd_sc_hd__buf_2 fanout147 (.A(net148),
    .X(net147));
 sky130_fd_sc_hd__buf_2 fanout148 (.A(\u_usb_host.u_core.fifo_rx_data_w[4] ),
    .X(net148));
 sky130_fd_sc_hd__buf_2 fanout149 (.A(net150),
    .X(net149));
 sky130_fd_sc_hd__buf_2 fanout150 (.A(\u_usb_host.u_core.fifo_rx_data_w[4] ),
    .X(net150));
 sky130_fd_sc_hd__buf_2 fanout151 (.A(net153),
    .X(net151));
 sky130_fd_sc_hd__buf_2 fanout152 (.A(net153),
    .X(net152));
 sky130_fd_sc_hd__buf_2 fanout153 (.A(net158),
    .X(net153));
 sky130_fd_sc_hd__buf_2 fanout154 (.A(net155),
    .X(net154));
 sky130_fd_sc_hd__buf_2 fanout155 (.A(net158),
    .X(net155));
 sky130_fd_sc_hd__buf_2 fanout156 (.A(net157),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 fanout157 (.A(net158),
    .X(net157));
 sky130_fd_sc_hd__clkbuf_4 fanout158 (.A(\u_usb_host.u_core.fifo_rx_data_w[3] ),
    .X(net158));
 sky130_fd_sc_hd__buf_2 fanout159 (.A(net161),
    .X(net159));
 sky130_fd_sc_hd__buf_2 fanout160 (.A(net161),
    .X(net160));
 sky130_fd_sc_hd__buf_2 fanout161 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net161));
 sky130_fd_sc_hd__buf_2 fanout162 (.A(net163),
    .X(net162));
 sky130_fd_sc_hd__buf_2 fanout163 (.A(net166),
    .X(net163));
 sky130_fd_sc_hd__buf_2 fanout164 (.A(net165),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_4 fanout165 (.A(net166),
    .X(net165));
 sky130_fd_sc_hd__clkbuf_2 fanout166 (.A(\u_usb_host.u_core.fifo_rx_data_w[2] ),
    .X(net166));
 sky130_fd_sc_hd__buf_2 fanout167 (.A(net168),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 fanout168 (.A(\u_usb_host.u_core.fifo_rx_data_w[1] ),
    .X(net168));
 sky130_fd_sc_hd__buf_2 fanout169 (.A(\u_usb_host.u_core.fifo_rx_data_w[1] ),
    .X(net169));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout170 (.A(\u_usb_host.u_core.fifo_rx_data_w[1] ),
    .X(net170));
 sky130_fd_sc_hd__buf_2 fanout171 (.A(net174),
    .X(net171));
 sky130_fd_sc_hd__buf_2 fanout172 (.A(net174),
    .X(net172));
 sky130_fd_sc_hd__buf_2 fanout173 (.A(net174),
    .X(net173));
 sky130_fd_sc_hd__buf_2 fanout174 (.A(\u_usb_host.u_core.fifo_rx_data_w[1] ),
    .X(net174));
 sky130_fd_sc_hd__buf_2 fanout175 (.A(net177),
    .X(net175));
 sky130_fd_sc_hd__buf_2 fanout176 (.A(net177),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_4 fanout177 (.A(\u_usb_host.u_core.fifo_rx_data_w[0] ),
    .X(net177));
 sky130_fd_sc_hd__buf_2 fanout178 (.A(net179),
    .X(net178));
 sky130_fd_sc_hd__buf_2 fanout179 (.A(net182),
    .X(net179));
 sky130_fd_sc_hd__buf_2 fanout180 (.A(net182),
    .X(net180));
 sky130_fd_sc_hd__clkbuf_2 fanout181 (.A(net182),
    .X(net181));
 sky130_fd_sc_hd__clkbuf_4 fanout182 (.A(\u_usb_host.u_core.fifo_rx_data_w[0] ),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_4 fanout183 (.A(\u_usb_host.u_core.u_sie._137_ ),
    .X(net183));
 sky130_fd_sc_hd__clkbuf_4 fanout184 (.A(\u_usb_host.u_core.u_fifo_tx._0575_ ),
    .X(net184));
 sky130_fd_sc_hd__clkbuf_2 fanout185 (.A(net187),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout186 (.A(net187),
    .X(net186));
 sky130_fd_sc_hd__clkbuf_4 fanout187 (.A(net188),
    .X(net187));
 sky130_fd_sc_hd__clkbuf_4 fanout188 (.A(\u_usb_host.u_core.u_fifo_tx._0573_ ),
    .X(net188));
 sky130_fd_sc_hd__buf_2 fanout189 (.A(net191),
    .X(net189));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout190 (.A(net191),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_4 fanout191 (.A(\u_usb_host.u_core.u_fifo_tx._0571_ ),
    .X(net191));
 sky130_fd_sc_hd__buf_2 fanout192 (.A(net193),
    .X(net192));
 sky130_fd_sc_hd__buf_2 fanout193 (.A(net194),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_2 fanout194 (.A(net195),
    .X(net194));
 sky130_fd_sc_hd__buf_2 fanout195 (.A(\u_usb_host.u_core.u_fifo_tx._0566_ ),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_2 fanout196 (.A(net197),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_2 fanout197 (.A(net198),
    .X(net197));
 sky130_fd_sc_hd__clkbuf_2 fanout198 (.A(net199),
    .X(net198));
 sky130_fd_sc_hd__buf_2 fanout199 (.A(\u_usb_host.u_core.u_fifo_tx._0563_ ),
    .X(net199));
 sky130_fd_sc_hd__clkbuf_2 fanout200 (.A(net201),
    .X(net200));
 sky130_fd_sc_hd__clkbuf_2 fanout201 (.A(net202),
    .X(net201));
 sky130_fd_sc_hd__buf_2 fanout202 (.A(\u_usb_host.u_core.u_fifo_tx._0549_ ),
    .X(net202));
 sky130_fd_sc_hd__clkbuf_2 fanout203 (.A(\u_usb_host.u_core.u_fifo_tx._0544_ ),
    .X(net203));
 sky130_fd_sc_hd__clkbuf_1 fanout204 (.A(\u_usb_host.u_core.u_fifo_tx._0544_ ),
    .X(net204));
 sky130_fd_sc_hd__clkbuf_2 fanout205 (.A(net206),
    .X(net205));
 sky130_fd_sc_hd__clkbuf_2 fanout206 (.A(net207),
    .X(net206));
 sky130_fd_sc_hd__clkbuf_4 fanout207 (.A(\u_usb_host.u_core.u_fifo_tx._0531_ ),
    .X(net207));
 sky130_fd_sc_hd__buf_2 fanout208 (.A(\u_usb_host.u_core.u_fifo_tx._0529_ ),
    .X(net208));
 sky130_fd_sc_hd__clkbuf_2 fanout209 (.A(\u_usb_host.u_core.u_fifo_tx._0529_ ),
    .X(net209));
 sky130_fd_sc_hd__clkbuf_4 fanout210 (.A(\u_usb_host.u_core.u_fifo_tx._0527_ ),
    .X(net210));
 sky130_fd_sc_hd__clkbuf_2 fanout211 (.A(net212),
    .X(net211));
 sky130_fd_sc_hd__clkbuf_2 fanout212 (.A(\u_usb_host.u_core.u_fifo_tx._0525_ ),
    .X(net212));
 sky130_fd_sc_hd__buf_2 fanout213 (.A(net215),
    .X(net213));
 sky130_fd_sc_hd__clkbuf_2 fanout214 (.A(net215),
    .X(net214));
 sky130_fd_sc_hd__buf_2 fanout215 (.A(net228),
    .X(net215));
 sky130_fd_sc_hd__clkbuf_2 fanout216 (.A(net218),
    .X(net216));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout217 (.A(net218),
    .X(net217));
 sky130_fd_sc_hd__clkbuf_2 fanout218 (.A(net219),
    .X(net218));
 sky130_fd_sc_hd__clkbuf_2 fanout219 (.A(net228),
    .X(net219));
 sky130_fd_sc_hd__clkbuf_2 fanout220 (.A(net221),
    .X(net220));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout221 (.A(net228),
    .X(net221));
 sky130_fd_sc_hd__clkbuf_2 fanout222 (.A(net228),
    .X(net222));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout223 (.A(net224),
    .X(net223));
 sky130_fd_sc_hd__clkbuf_2 fanout224 (.A(net228),
    .X(net224));
 sky130_fd_sc_hd__clkbuf_2 fanout225 (.A(net227),
    .X(net225));
 sky130_fd_sc_hd__clkbuf_1 fanout226 (.A(net227),
    .X(net226));
 sky130_fd_sc_hd__clkbuf_2 fanout227 (.A(net228),
    .X(net227));
 sky130_fd_sc_hd__clkbuf_4 fanout228 (.A(\u_usb_host.u_core.u_fifo_tx._0523_ ),
    .X(net228));
 sky130_fd_sc_hd__clkbuf_4 fanout229 (.A(net231),
    .X(net229));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout230 (.A(net231),
    .X(net230));
 sky130_fd_sc_hd__clkbuf_4 fanout231 (.A(\u_usb_host.u_core.u_fifo_tx._0522_ ),
    .X(net231));
 sky130_fd_sc_hd__buf_2 fanout232 (.A(\u_usb_host.u_core.u_fifo_tx._0520_ ),
    .X(net232));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout233 (.A(\u_usb_host.u_core.u_fifo_tx._0520_ ),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_2 fanout234 (.A(net235),
    .X(net234));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout235 (.A(net238),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_2 fanout236 (.A(net238),
    .X(net236));
 sky130_fd_sc_hd__buf_2 fanout237 (.A(net238),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_2 fanout238 (.A(net240),
    .X(net238));
 sky130_fd_sc_hd__buf_2 fanout239 (.A(net240),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_2 fanout240 (.A(\u_usb_host.u_core.u_fifo_tx._0517_ ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_2 fanout241 (.A(net243),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 fanout242 (.A(net243),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_4 fanout243 (.A(\u_usb_host.u_core.u_fifo_tx._0516_ ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_2 fanout244 (.A(net258),
    .X(net244));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout245 (.A(net258),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_2 fanout246 (.A(net247),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_2 fanout247 (.A(net250),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_2 fanout248 (.A(net249),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_2 fanout249 (.A(net250),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_2 fanout250 (.A(net258),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_2 fanout251 (.A(net256),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 fanout252 (.A(net256),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_2 fanout253 (.A(net255),
    .X(net253));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout254 (.A(net255),
    .X(net254));
 sky130_fd_sc_hd__clkbuf_2 fanout255 (.A(net256),
    .X(net255));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout256 (.A(net257),
    .X(net256));
 sky130_fd_sc_hd__clkbuf_2 fanout257 (.A(net258),
    .X(net257));
 sky130_fd_sc_hd__clkbuf_4 fanout258 (.A(\u_usb_host.u_core.u_fifo_tx._0509_ ),
    .X(net258));
 sky130_fd_sc_hd__clkbuf_2 fanout259 (.A(net261),
    .X(net259));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout260 (.A(net261),
    .X(net260));
 sky130_fd_sc_hd__buf_2 fanout261 (.A(\u_usb_host.u_core.u_fifo_tx._0508_ ),
    .X(net261));
 sky130_fd_sc_hd__clkbuf_2 fanout262 (.A(net264),
    .X(net262));
 sky130_fd_sc_hd__clkbuf_2 fanout263 (.A(net264),
    .X(net263));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout264 (.A(net266),
    .X(net264));
 sky130_fd_sc_hd__clkbuf_2 fanout265 (.A(net266),
    .X(net265));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout266 (.A(\u_usb_host.u_core.u_fifo_tx._0508_ ),
    .X(net266));
 sky130_fd_sc_hd__clkbuf_2 fanout267 (.A(net268),
    .X(net267));
 sky130_fd_sc_hd__buf_2 fanout268 (.A(\u_usb_host.u_core.u_fifo_tx._0508_ ),
    .X(net268));
 sky130_fd_sc_hd__buf_2 fanout269 (.A(net270),
    .X(net269));
 sky130_fd_sc_hd__buf_2 fanout270 (.A(net273),
    .X(net270));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout271 (.A(net273),
    .X(net271));
 sky130_fd_sc_hd__clkbuf_2 fanout272 (.A(net273),
    .X(net272));
 sky130_fd_sc_hd__buf_2 fanout273 (.A(\u_usb_host.u_core.u_fifo_tx._0506_ ),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_4 fanout274 (.A(\u_usb_host.u_core.u_fifo_tx._0504_ ),
    .X(net274));
 sky130_fd_sc_hd__buf_2 fanout275 (.A(\u_usb_host.u_core.u_fifo_rx._0575_ ),
    .X(net275));
 sky130_fd_sc_hd__clkbuf_2 fanout276 (.A(\u_usb_host.u_core.u_fifo_rx._0573_ ),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 fanout277 (.A(\u_usb_host.u_core.u_fifo_rx._0573_ ),
    .X(net277));
 sky130_fd_sc_hd__buf_2 fanout278 (.A(net279),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_2 fanout279 (.A(\u_usb_host.u_core.u_fifo_rx._0573_ ),
    .X(net279));
 sky130_fd_sc_hd__buf_2 fanout280 (.A(net282),
    .X(net280));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout281 (.A(net282),
    .X(net281));
 sky130_fd_sc_hd__clkbuf_4 fanout282 (.A(\u_usb_host.u_core.u_fifo_rx._0571_ ),
    .X(net282));
 sky130_fd_sc_hd__clkbuf_2 fanout283 (.A(\u_usb_host.u_core.u_fifo_rx._0566_ ),
    .X(net283));
 sky130_fd_sc_hd__clkbuf_1 fanout284 (.A(\u_usb_host.u_core.u_fifo_rx._0566_ ),
    .X(net284));
 sky130_fd_sc_hd__buf_2 fanout285 (.A(\u_usb_host.u_core.u_fifo_rx._0566_ ),
    .X(net285));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout286 (.A(\u_usb_host.u_core.u_fifo_rx._0566_ ),
    .X(net286));
 sky130_fd_sc_hd__clkbuf_4 fanout287 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net287));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout288 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net288));
 sky130_fd_sc_hd__buf_2 fanout289 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net289));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout290 (.A(\u_usb_host.u_core.u_fifo_rx._0563_ ),
    .X(net290));
 sky130_fd_sc_hd__clkbuf_2 fanout291 (.A(net292),
    .X(net291));
 sky130_fd_sc_hd__clkbuf_2 fanout292 (.A(net293),
    .X(net292));
 sky130_fd_sc_hd__clkbuf_4 fanout293 (.A(\u_usb_host.u_core.u_fifo_rx._0549_ ),
    .X(net293));
 sky130_fd_sc_hd__buf_2 fanout294 (.A(\u_usb_host.u_core.u_fifo_rx._0544_ ),
    .X(net294));
 sky130_fd_sc_hd__buf_2 fanout295 (.A(\u_usb_host.u_core.u_fifo_rx._0544_ ),
    .X(net295));
 sky130_fd_sc_hd__buf_2 fanout296 (.A(net298),
    .X(net296));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout297 (.A(net298),
    .X(net297));
 sky130_fd_sc_hd__buf_4 fanout298 (.A(\u_usb_host.u_core.u_fifo_rx._0531_ ),
    .X(net298));
 sky130_fd_sc_hd__clkbuf_4 fanout299 (.A(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .X(net299));
 sky130_fd_sc_hd__clkbuf_2 fanout300 (.A(\u_usb_host.u_core.u_fifo_rx._0529_ ),
    .X(net300));
 sky130_fd_sc_hd__clkbuf_4 fanout301 (.A(\u_usb_host.u_core.u_fifo_rx._0527_ ),
    .X(net301));
 sky130_fd_sc_hd__clkbuf_2 fanout302 (.A(net303),
    .X(net302));
 sky130_fd_sc_hd__clkbuf_2 fanout303 (.A(\u_usb_host.u_core.u_fifo_rx._0525_ ),
    .X(net303));
 sky130_fd_sc_hd__clkbuf_2 fanout304 (.A(net305),
    .X(net304));
 sky130_fd_sc_hd__clkbuf_2 fanout305 (.A(net306),
    .X(net305));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout306 (.A(net310),
    .X(net306));
 sky130_fd_sc_hd__clkbuf_2 fanout307 (.A(net308),
    .X(net307));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout308 (.A(net309),
    .X(net308));
 sky130_fd_sc_hd__clkbuf_2 fanout309 (.A(net310),
    .X(net309));
 sky130_fd_sc_hd__clkbuf_2 fanout310 (.A(\u_usb_host.u_core.u_fifo_rx._0523_ ),
    .X(net310));
 sky130_fd_sc_hd__clkbuf_2 fanout311 (.A(net312),
    .X(net311));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout312 (.A(net319),
    .X(net312));
 sky130_fd_sc_hd__clkbuf_2 fanout313 (.A(net318),
    .X(net313));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout314 (.A(net318),
    .X(net314));
 sky130_fd_sc_hd__clkbuf_2 fanout315 (.A(net318),
    .X(net315));
 sky130_fd_sc_hd__clkbuf_2 fanout316 (.A(net317),
    .X(net316));
 sky130_fd_sc_hd__clkbuf_2 fanout317 (.A(net318),
    .X(net317));
 sky130_fd_sc_hd__clkbuf_2 fanout318 (.A(net319),
    .X(net318));
 sky130_fd_sc_hd__buf_2 fanout319 (.A(\u_usb_host.u_core.u_fifo_rx._0523_ ),
    .X(net319));
 sky130_fd_sc_hd__buf_2 fanout320 (.A(net322),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 fanout321 (.A(net322),
    .X(net321));
 sky130_fd_sc_hd__buf_2 fanout322 (.A(\u_usb_host.u_core.u_fifo_rx._0522_ ),
    .X(net322));
 sky130_fd_sc_hd__clkbuf_4 fanout323 (.A(\u_usb_host.u_core.u_fifo_rx._0520_ ),
    .X(net323));
 sky130_fd_sc_hd__clkbuf_2 fanout324 (.A(\u_usb_host.u_core.u_fifo_rx._0520_ ),
    .X(net324));
 sky130_fd_sc_hd__clkbuf_2 fanout325 (.A(net327),
    .X(net325));
 sky130_fd_sc_hd__clkbuf_1 fanout326 (.A(net327),
    .X(net326));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout327 (.A(net328),
    .X(net327));
 sky130_fd_sc_hd__clkbuf_2 fanout328 (.A(net329),
    .X(net328));
 sky130_fd_sc_hd__buf_2 fanout329 (.A(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .X(net329));
 sky130_fd_sc_hd__buf_2 fanout330 (.A(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .X(net330));
 sky130_fd_sc_hd__clkbuf_1 fanout331 (.A(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_2 fanout332 (.A(net333),
    .X(net332));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout333 (.A(net334),
    .X(net333));
 sky130_fd_sc_hd__clkbuf_4 fanout334 (.A(\u_usb_host.u_core.u_fifo_rx._0516_ ),
    .X(net334));
 sky130_fd_sc_hd__clkbuf_2 fanout335 (.A(net337),
    .X(net335));
 sky130_fd_sc_hd__clkbuf_1 fanout336 (.A(net337),
    .X(net336));
 sky130_fd_sc_hd__buf_2 fanout337 (.A(\u_usb_host.u_core.u_fifo_rx._0509_ ),
    .X(net337));
 sky130_fd_sc_hd__clkbuf_2 fanout338 (.A(net348),
    .X(net338));
 sky130_fd_sc_hd__clkbuf_2 fanout339 (.A(net341),
    .X(net339));
 sky130_fd_sc_hd__clkbuf_2 fanout340 (.A(net341),
    .X(net340));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout341 (.A(net348),
    .X(net341));
 sky130_fd_sc_hd__clkbuf_2 fanout342 (.A(net347),
    .X(net342));
 sky130_fd_sc_hd__clkbuf_2 fanout343 (.A(net346),
    .X(net343));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout344 (.A(net346),
    .X(net344));
 sky130_fd_sc_hd__clkbuf_2 fanout345 (.A(net346),
    .X(net345));
 sky130_fd_sc_hd__clkbuf_2 fanout346 (.A(net347),
    .X(net346));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout347 (.A(net348),
    .X(net347));
 sky130_fd_sc_hd__buf_2 fanout348 (.A(\u_usb_host.u_core.u_fifo_rx._0509_ ),
    .X(net348));
 sky130_fd_sc_hd__clkbuf_2 fanout349 (.A(net350),
    .X(net349));
 sky130_fd_sc_hd__clkbuf_2 fanout350 (.A(net352),
    .X(net350));
 sky130_fd_sc_hd__clkbuf_2 fanout351 (.A(net352),
    .X(net351));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout352 (.A(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .X(net352));
 sky130_fd_sc_hd__clkbuf_2 fanout353 (.A(net354),
    .X(net353));
 sky130_fd_sc_hd__clkbuf_2 fanout354 (.A(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .X(net354));
 sky130_fd_sc_hd__clkbuf_2 fanout355 (.A(net358),
    .X(net355));
 sky130_fd_sc_hd__clkbuf_2 fanout356 (.A(net358),
    .X(net356));
 sky130_fd_sc_hd__buf_2 fanout357 (.A(net358),
    .X(net357));
 sky130_fd_sc_hd__clkbuf_2 fanout358 (.A(\u_usb_host.u_core.u_fifo_rx._0508_ ),
    .X(net358));
 sky130_fd_sc_hd__clkbuf_2 fanout359 (.A(net361),
    .X(net359));
 sky130_fd_sc_hd__clkbuf_2 fanout360 (.A(net361),
    .X(net360));
 sky130_fd_sc_hd__clkbuf_2 fanout361 (.A(\u_usb_host.u_core.u_fifo_rx._0506_ ),
    .X(net361));
 sky130_fd_sc_hd__buf_2 fanout362 (.A(\u_usb_host.u_core.u_fifo_rx._0506_ ),
    .X(net362));
 sky130_fd_sc_hd__buf_4 fanout363 (.A(\u_usb_host.u_core.u_fifo_rx._0504_ ),
    .X(net363));
 sky130_fd_sc_hd__clkbuf_4 fanout364 (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .X(net364));
 sky130_fd_sc_hd__clkbuf_4 fanout365 (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .X(net365));
 sky130_fd_sc_hd__clkbuf_4 fanout366 (.A(net367),
    .X(net366));
 sky130_fd_sc_hd__clkbuf_4 fanout367 (.A(net372),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_4 fanout368 (.A(net372),
    .X(net368));
 sky130_fd_sc_hd__clkbuf_4 fanout369 (.A(net372),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_4 fanout370 (.A(net371),
    .X(net370));
 sky130_fd_sc_hd__buf_2 fanout371 (.A(net372),
    .X(net371));
 sky130_fd_sc_hd__buf_2 fanout372 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_4 fanout373 (.A(net374),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 fanout374 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_4 fanout375 (.A(net376),
    .X(net375));
 sky130_fd_sc_hd__buf_2 fanout376 (.A(net377),
    .X(net376));
 sky130_fd_sc_hd__buf_2 fanout377 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_4 fanout378 (.A(net379),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_2 fanout379 (.A(net386),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_4 fanout380 (.A(net381),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_2 fanout381 (.A(net386),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_4 fanout382 (.A(net386),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_4 fanout383 (.A(net386),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_4 fanout384 (.A(net386),
    .X(net384));
 sky130_fd_sc_hd__clkbuf_2 fanout385 (.A(net386),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_2 fanout386 (.A(net416),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_4 fanout387 (.A(net388),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_4 fanout388 (.A(net392),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_4 fanout389 (.A(net392),
    .X(net389));
 sky130_fd_sc_hd__buf_2 fanout390 (.A(net392),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_4 fanout391 (.A(net392),
    .X(net391));
 sky130_fd_sc_hd__buf_2 fanout392 (.A(net416),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_4 fanout393 (.A(net395),
    .X(net393));
 sky130_fd_sc_hd__buf_2 fanout394 (.A(net395),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_4 fanout395 (.A(net416),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_4 fanout396 (.A(net397),
    .X(net396));
 sky130_fd_sc_hd__buf_2 fanout397 (.A(net398),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_4 fanout398 (.A(net403),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_4 fanout399 (.A(net400),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_4 fanout400 (.A(net403),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_4 fanout401 (.A(net402),
    .X(net401));
 sky130_fd_sc_hd__buf_2 fanout402 (.A(net403),
    .X(net402));
 sky130_fd_sc_hd__buf_2 fanout403 (.A(net416),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_4 fanout404 (.A(net415),
    .X(net404));
 sky130_fd_sc_hd__buf_2 fanout405 (.A(net415),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_4 fanout406 (.A(net409),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_4 fanout407 (.A(net408),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_4 fanout408 (.A(net409),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_2 fanout409 (.A(net415),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_4 fanout410 (.A(net411),
    .X(net410));
 sky130_fd_sc_hd__buf_2 fanout411 (.A(net415),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_4 fanout412 (.A(net413),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_4 fanout413 (.A(net414),
    .X(net413));
 sky130_fd_sc_hd__buf_2 fanout414 (.A(net415),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_2 fanout415 (.A(net416),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_4 fanout416 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ),
    .X(net416));
 sky130_fd_sc_hd__buf_2 fanout417 (.A(\u_usb_host.u_phy.state_q[3] ),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_2 fanout418 (.A(\u_usb_host.u_phy.state_q[2] ),
    .X(net418));
 sky130_fd_sc_hd__buf_2 fanout419 (.A(\u_usb_host.u_phy.state_q[1] ),
    .X(net419));
 sky130_fd_sc_hd__clkbuf_1 fanout420 (.A(\u_usb_host.u_phy.state_q[1] ),
    .X(net420));
 sky130_fd_sc_hd__buf_2 fanout421 (.A(\u_usb_host.u_phy.state_q[0] ),
    .X(net421));
 sky130_fd_sc_hd__buf_2 fanout422 (.A(net424),
    .X(net422));
 sky130_fd_sc_hd__buf_2 fanout423 (.A(net424),
    .X(net423));
 sky130_fd_sc_hd__buf_2 fanout424 (.A(\u_usb_host.u_core.u_sie._120_ ),
    .X(net424));
 sky130_fd_sc_hd__buf_4 fanout425 (.A(\u_usb_host.u_core.u_sie._082_ ),
    .X(net425));
 sky130_fd_sc_hd__buf_2 fanout426 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[3] ),
    .X(net426));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout427 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[3] ),
    .X(net427));
 sky130_fd_sc_hd__clkbuf_2 fanout428 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ),
    .X(net428));
 sky130_fd_sc_hd__buf_2 fanout429 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[1] ),
    .X(net429));
 sky130_fd_sc_hd__clkbuf_2 fanout430 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[1] ),
    .X(net430));
 sky130_fd_sc_hd__clkbuf_2 fanout431 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[0] ),
    .X(net431));
 sky130_fd_sc_hd__buf_2 fanout432 (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[0] ),
    .X(net432));
 sky130_fd_sc_hd__buf_2 fanout433 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[3] ),
    .X(net433));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout434 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[3] ),
    .X(net434));
 sky130_fd_sc_hd__buf_2 fanout435 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[2] ),
    .X(net435));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout436 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[2] ),
    .X(net436));
 sky130_fd_sc_hd__clkbuf_2 fanout437 (.A(net438),
    .X(net437));
 sky130_fd_sc_hd__clkbuf_4 fanout438 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[1] ),
    .X(net438));
 sky130_fd_sc_hd__clkbuf_2 fanout439 (.A(net440),
    .X(net439));
 sky130_fd_sc_hd__clkbuf_4 fanout440 (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[0] ),
    .X(net440));
 sky130_fd_sc_hd__buf_2 fanout441 (.A(net442),
    .X(net441));
 sky130_fd_sc_hd__clkbuf_2 fanout442 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ),
    .X(net442));
 sky130_fd_sc_hd__clkbuf_2 fanout443 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .X(net443));
 sky130_fd_sc_hd__clkbuf_2 fanout444 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .X(net444));
 sky130_fd_sc_hd__clkbuf_2 fanout445 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ),
    .X(net445));
 sky130_fd_sc_hd__buf_2 fanout446 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .X(net446));
 sky130_fd_sc_hd__clkbuf_2 fanout447 (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ),
    .X(net447));
 sky130_fd_sc_hd__buf_2 fanout448 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ),
    .X(net448));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout449 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ),
    .X(net449));
 sky130_fd_sc_hd__buf_2 fanout450 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ),
    .X(net450));
 sky130_fd_sc_hd__buf_2 fanout451 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ),
    .X(net451));
 sky130_fd_sc_hd__buf_2 fanout452 (.A(net453),
    .X(net452));
 sky130_fd_sc_hd__clkbuf_2 fanout453 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ),
    .X(net453));
 sky130_fd_sc_hd__buf_2 fanout454 (.A(net456),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_2 fanout455 (.A(net456),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_2 fanout456 (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ),
    .X(net456));
 sky130_fd_sc_hd__buf_2 fanout457 (.A(net465),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_2 fanout458 (.A(net465),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_4 fanout459 (.A(net465),
    .X(net459));
 sky130_fd_sc_hd__clkbuf_2 fanout460 (.A(net465),
    .X(net460));
 sky130_fd_sc_hd__clkbuf_4 fanout461 (.A(net464),
    .X(net461));
 sky130_fd_sc_hd__buf_2 fanout462 (.A(net464),
    .X(net462));
 sky130_fd_sc_hd__buf_2 fanout463 (.A(net464),
    .X(net463));
 sky130_fd_sc_hd__clkbuf_2 fanout464 (.A(net465),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_4 fanout465 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[7] ),
    .X(net465));
 sky130_fd_sc_hd__clkbuf_4 fanout466 (.A(net473),
    .X(net466));
 sky130_fd_sc_hd__clkbuf_2 fanout467 (.A(net473),
    .X(net467));
 sky130_fd_sc_hd__buf_2 fanout468 (.A(net473),
    .X(net468));
 sky130_fd_sc_hd__buf_2 fanout469 (.A(net473),
    .X(net469));
 sky130_fd_sc_hd__buf_2 fanout470 (.A(net471),
    .X(net470));
 sky130_fd_sc_hd__buf_2 fanout471 (.A(net472),
    .X(net471));
 sky130_fd_sc_hd__clkbuf_4 fanout472 (.A(net473),
    .X(net472));
 sky130_fd_sc_hd__buf_4 fanout473 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[6] ),
    .X(net473));
 sky130_fd_sc_hd__clkbuf_4 fanout474 (.A(net482),
    .X(net474));
 sky130_fd_sc_hd__clkbuf_2 fanout475 (.A(net482),
    .X(net475));
 sky130_fd_sc_hd__clkbuf_4 fanout476 (.A(net482),
    .X(net476));
 sky130_fd_sc_hd__clkbuf_2 fanout477 (.A(net482),
    .X(net477));
 sky130_fd_sc_hd__clkbuf_4 fanout478 (.A(net481),
    .X(net478));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout479 (.A(net481),
    .X(net479));
 sky130_fd_sc_hd__buf_2 fanout480 (.A(net481),
    .X(net480));
 sky130_fd_sc_hd__buf_2 fanout481 (.A(net482),
    .X(net481));
 sky130_fd_sc_hd__clkbuf_4 fanout482 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[5] ),
    .X(net482));
 sky130_fd_sc_hd__buf_2 fanout483 (.A(net484),
    .X(net483));
 sky130_fd_sc_hd__clkbuf_4 fanout484 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[4] ),
    .X(net484));
 sky130_fd_sc_hd__clkbuf_4 fanout485 (.A(net486),
    .X(net485));
 sky130_fd_sc_hd__clkbuf_4 fanout486 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[4] ),
    .X(net486));
 sky130_fd_sc_hd__clkbuf_4 fanout487 (.A(net490),
    .X(net487));
 sky130_fd_sc_hd__clkbuf_2 fanout488 (.A(net490),
    .X(net488));
 sky130_fd_sc_hd__clkbuf_4 fanout489 (.A(net490),
    .X(net489));
 sky130_fd_sc_hd__buf_2 fanout490 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[4] ),
    .X(net490));
 sky130_fd_sc_hd__clkbuf_4 fanout491 (.A(net499),
    .X(net491));
 sky130_fd_sc_hd__clkbuf_2 fanout492 (.A(net499),
    .X(net492));
 sky130_fd_sc_hd__clkbuf_4 fanout493 (.A(net499),
    .X(net493));
 sky130_fd_sc_hd__buf_2 fanout494 (.A(net499),
    .X(net494));
 sky130_fd_sc_hd__clkbuf_4 fanout495 (.A(net498),
    .X(net495));
 sky130_fd_sc_hd__buf_2 fanout496 (.A(net498),
    .X(net496));
 sky130_fd_sc_hd__buf_2 fanout497 (.A(net498),
    .X(net497));
 sky130_fd_sc_hd__buf_2 fanout498 (.A(net499),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_4 fanout499 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[3] ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_4 fanout500 (.A(net508),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_2 fanout501 (.A(net508),
    .X(net501));
 sky130_fd_sc_hd__clkbuf_4 fanout502 (.A(net508),
    .X(net502));
 sky130_fd_sc_hd__buf_2 fanout503 (.A(net508),
    .X(net503));
 sky130_fd_sc_hd__clkbuf_4 fanout504 (.A(net508),
    .X(net504));
 sky130_fd_sc_hd__clkbuf_2 fanout505 (.A(net508),
    .X(net505));
 sky130_fd_sc_hd__clkbuf_4 fanout506 (.A(net507),
    .X(net506));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout507 (.A(net508),
    .X(net507));
 sky130_fd_sc_hd__buf_4 fanout508 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[2] ),
    .X(net508));
 sky130_fd_sc_hd__buf_2 fanout509 (.A(net510),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_2 fanout510 (.A(net513),
    .X(net510));
 sky130_fd_sc_hd__buf_2 fanout511 (.A(net513),
    .X(net511));
 sky130_fd_sc_hd__buf_2 fanout512 (.A(net513),
    .X(net512));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[1] ),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_4 fanout514 (.A(net516),
    .X(net514));
 sky130_fd_sc_hd__buf_2 fanout515 (.A(net516),
    .X(net515));
 sky130_fd_sc_hd__clkbuf_4 fanout516 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[1] ),
    .X(net516));
 sky130_fd_sc_hd__buf_2 fanout517 (.A(net520),
    .X(net517));
 sky130_fd_sc_hd__buf_2 fanout518 (.A(net519),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_4 fanout519 (.A(net520),
    .X(net519));
 sky130_fd_sc_hd__buf_4 fanout520 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[0] ),
    .X(net520));
 sky130_fd_sc_hd__buf_2 fanout521 (.A(net522),
    .X(net521));
 sky130_fd_sc_hd__clkbuf_4 fanout522 (.A(net523),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_4 fanout523 (.A(\u_usb_host.u_core.u_fifo_tx.data_i[0] ),
    .X(net523));
 sky130_fd_sc_hd__clkbuf_4 fanout524 (.A(net525),
    .X(net524));
 sky130_fd_sc_hd__buf_2 fanout525 (.A(\u_usb_host.u_core.sof_transfer_q ),
    .X(net525));
 sky130_fd_sc_hd__clkbuf_4 fanout526 (.A(net569),
    .X(net526));
 sky130_fd_sc_hd__buf_2 fanout527 (.A(net569),
    .X(net527));
 sky130_fd_sc_hd__clkbuf_4 fanout528 (.A(net569),
    .X(net528));
 sky130_fd_sc_hd__buf_2 fanout529 (.A(net568),
    .X(net529));
 sky130_fd_sc_hd__buf_2 fanout530 (.A(net567),
    .X(net530));
 sky130_fd_sc_hd__clkbuf_4 fanout531 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ),
    .X(net531));
 sky130_fd_sc_hd__clkbuf_4 fanout532 (.A(net534),
    .X(net532));
 sky130_fd_sc_hd__clkbuf_4 fanout533 (.A(net534),
    .X(net533));
 sky130_fd_sc_hd__clkbuf_4 fanout534 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ),
    .X(net534));
 sky130_fd_sc_hd__buf_4 fanout535 (.A(net539),
    .X(net535));
 sky130_fd_sc_hd__buf_4 fanout536 (.A(net538),
    .X(net536));
 sky130_fd_sc_hd__buf_4 fanout537 (.A(net538),
    .X(net537));
 sky130_fd_sc_hd__buf_4 fanout538 (.A(net539),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_2 fanout539 (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(\u_usb_host.u_core.u_sie.utmi_txready_i ),
    .X(net540));
 sky130_fd_sc_hd__buf_2 fanout541 (.A(net542),
    .X(net541));
 sky130_fd_sc_hd__clkbuf_2 fanout542 (.A(\u_usb_host.u_core.u_sie.state_q[1] ),
    .X(net542));
 sky130_fd_sc_hd__buf_2 fanout543 (.A(\u_usb_host.u_core.u_sie.state_q[0] ),
    .X(net543));
 sky130_fd_sc_hd__buf_2 fanout86 (.A(net87),
    .X(net86));
 sky130_fd_sc_hd__buf_2 fanout87 (.A(net88),
    .X(net87));
 sky130_fd_sc_hd__clkbuf_4 fanout88 (.A(\u_usb_host.u_core._117_ ),
    .X(net88));
 sky130_fd_sc_hd__buf_2 fanout89 (.A(net91),
    .X(net89));
 sky130_fd_sc_hd__clkbuf_2 fanout90 (.A(net91),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_2 fanout91 (.A(\u_usb_host.u_core._099_ ),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_4 fanout92 (.A(\u_usb_host.u_core._097_ ),
    .X(net92));
 sky130_fd_sc_hd__buf_2 fanout93 (.A(\u_usb_host.u_core._097_ ),
    .X(net93));
 sky130_fd_sc_hd__buf_2 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__clkbuf_2 fanout95 (.A(net96),
    .X(net95));
 sky130_fd_sc_hd__buf_2 fanout96 (.A(\u_usb_host.u_core._091_ ),
    .X(net96));
 sky130_fd_sc_hd__buf_4 fanout97 (.A(\u_usb_host.u_core.u_fifo_rx._0475_ ),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 fanout98 (.A(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .X(net98));
 sky130_fd_sc_hd__clkbuf_4 fanout99 (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ),
    .X(net567));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\u_usb_host.u_core.status_crc_err_w ),
    .X(net576));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[25] ),
    .X(net666));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[16] ),
    .X(net667));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\u_usb_host.reg_rdata[25] ),
    .X(net668));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[30] ),
    .X(net669));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[29] ),
    .X(net670));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\u_usb_host.u_phy.rxd_last_j_q ),
    .X(net671));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[14] ),
    .X(net672));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ),
    .X(net673));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ),
    .X(net674));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(\u_usb_host.u_core.u_sie.rx_active_q[1] ),
    .X(net675));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\u_usb_host.u_core.reg_rdata_r[30] ),
    .X(net577));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(\u_usb_host.u_core.u_sie.rx_active_q[2] ),
    .X(net676));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ),
    .X(net677));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\u_usb_host.u_phy.rxd_ms ),
    .X(net678));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ),
    .X(net679));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ),
    .X(net680));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ),
    .X(net681));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\u_usb_host.u_core.transfer_start_q ),
    .X(net682));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\u_usb_host.u_phy.rx_dp_ms ),
    .X(net683));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\u_usb_host.u_core.in_transfer_q ),
    .X(net684));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\u_usb_host.u_phy.rxd1_q ),
    .X(net685));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_usb_host.u_core.status_timeout_w ),
    .X(net578));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\u_usb_host.u_phy.rx_dp1_q ),
    .X(net686));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\u_usb_host.u_core.u_sie.data_ready_w ),
    .X(net687));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\u_usb_host.u_core.u_sie.data_idx_i ),
    .X(net688));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\u_usb_host.u_core.reg_rdata_r[29] ),
    .X(net579));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\u_usb_host.u_phy.rxd_last_q ),
    .X(net580));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u_usb_host.u_core.u_sie.se0_detect_q ),
    .X(net581));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\u_usb_host.u_core.u_sie._171_ ),
    .X(net582));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .X(net583));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u_usb_host.u_core.u_sie.utmi_txready_i ),
    .X(net584));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\u_usb_host.u_core.usb_err_q ),
    .X(net585));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(net530),
    .X(net568));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\u_usb_host.u_core.reg_rdata_r[2] ),
    .X(net586));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\u_usb_host.u_core.sof_irq_q ),
    .X(net587));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\u_usb_host.u_core.u_sie.data_idx_i ),
    .X(net588));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ),
    .X(net589));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u_usb_host.u_core.intr_done_q ),
    .X(net590));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\u_usb_host.u_core.reg_rdata_r[1] ),
    .X(net591));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\u_usb_host.u_core.usb_irq_mask_sof_out_w ),
    .X(net592));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\u_usb_host.u_core._131_ ),
    .X(net593));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\u_usb_host.u_core.utmi_termselect_o ),
    .X(net594));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\u_usb_host.u_phy.sync_j_detected_q ),
    .X(net595));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(net529),
    .X(net569));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_usb_host.reg_rdata[8] ),
    .X(net596));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\u_usb_host.reg_rdata[21] ),
    .X(net597));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\u_usb_host.reg_rdata[16] ),
    .X(net598));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\u_usb_host.reg_rdata[11] ),
    .X(net599));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\u_usb_host.reg_rdata[28] ),
    .X(net600));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\u_usb_host.u_core.utmi_dmpulldown_o ),
    .X(net601));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\u_usb_host.reg_rdata[22] ),
    .X(net602));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\u_usb_host.reg_rdata[13] ),
    .X(net603));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\u_usb_host.reg_rdata[9] ),
    .X(net604));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u_usb_host.reg_rdata[1] ),
    .X(net605));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net572),
    .X(net570));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\u_usb_host.reg_rdata[12] ),
    .X(net606));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\u_usb_host.reg_rdata[6] ),
    .X(net607));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u_usb_host.reg_rdata[0] ),
    .X(net608));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\u_usb_host.reg_rdata[2] ),
    .X(net609));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\u_usb_host.reg_rdata[31] ),
    .X(net610));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[3] ),
    .X(net611));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\u_usb_host.u_core.utmi_dppulldown_o ),
    .X(net612));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\u_usb_host.reg_rdata[29] ),
    .X(net613));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u_usb_host.u_core.usb_ctrl_wr_q ),
    .X(net614));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[7] ),
    .X(net615));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ),
    .X(net571));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[2] ),
    .X(net616));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u_usb_host.reg_rdata[5] ),
    .X(net617));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\u_usb_host.reg_rdata[3] ),
    .X(net618));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\u_usb_host.reg_rdata[7] ),
    .X(net619));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[4] ),
    .X(net620));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[5] ),
    .X(net621));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[1] ),
    .X(net622));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\u_usb_host.reg_rdata[4] ),
    .X(net623));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\u_usb_host.u_core.u_sie.utmi_data_i[6] ),
    .X(net624));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\u_usb_host.reg_rdata[18] ),
    .X(net625));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\u_usb_host.u_wb_rst.in_data_2s ),
    .X(net572));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\u_usb_host.reg_rdata[10] ),
    .X(net626));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\u_usb_host.reg_rdata[14] ),
    .X(net627));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\u_usb_host.reg_rdata[20] ),
    .X(net628));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\u_usb_host.reg_rdata[15] ),
    .X(net629));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\u_usb_host.reg_rdata[19] ),
    .X(net630));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\u_usb_host.u_core.u_sie.data_valid_q[3] ),
    .X(net631));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\u_usb_host.reg_rdata[27] ),
    .X(net632));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[19] ),
    .X(net633));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[17] ),
    .X(net634));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[21] ),
    .X(net635));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\u_usb_host.u_usb_rst.in_data_2s ),
    .X(net573));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[23] ),
    .X(net636));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[8] ),
    .X(net637));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[18] ),
    .X(net638));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[10] ),
    .X(net639));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(\u_usb_host.reg_rdata[30] ),
    .X(net640));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(\u_usb_host.u_core.u_sie.data_crc_q[1] ),
    .X(net641));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[20] ),
    .X(net642));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\u_usb_host.reg_rdata[26] ),
    .X(net643));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(\u_usb_host.reg_rdata[23] ),
    .X(net644));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(\u_usb_host.reg_rdata[17] ),
    .X(net645));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\u_usb_host.u_core.u_sie.utmi_rxvalid_i ),
    .X(net574));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(\u_usb_host.reg_rdata[24] ),
    .X(net646));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\u_usb_host.u_phy.rx_dn_ms ),
    .X(net647));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(\u_usb_host.u_usb_rst.in_data_s ),
    .X(net648));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[22] ),
    .X(net649));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[13] ),
    .X(net650));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[9] ),
    .X(net651));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[12] ),
    .X(net652));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[11] ),
    .X(net653));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[28] ),
    .X(net654));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ),
    .X(net655));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\u_usb_host.u_core.u_fifo_tx.push_i ),
    .X(net575));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ),
    .X(net656));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ),
    .X(net657));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ),
    .X(net658));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(\u_usb_host.u_wb_rst.in_data_s ),
    .X(net659));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(\u_usb_host.u_core.u_sie.data_valid_q[2] ),
    .X(net660));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[26] ),
    .X(net661));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[31] ),
    .X(net662));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[24] ),
    .X(net663));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[27] ),
    .X(net664));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\u_usb_host.u_core.u_sie.data_buffer_q[15] ),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 input1 (.A(cfg_cska_usb[0]),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(reg_addr[5]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(reg_addr[6]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(reg_addr[7]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(reg_addr[8]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(reg_cs),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_1 input15 (.A(reg_wdata[0]),
    .X(net15));
 sky130_fd_sc_hd__dlymetal6s2s_1 input16 (.A(reg_wdata[10]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(reg_wdata[11]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(reg_wdata[12]),
    .X(net18));
 sky130_fd_sc_hd__dlymetal6s2s_1 input19 (.A(reg_wdata[13]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(cfg_cska_usb[1]),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(reg_wdata[14]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_1 input21 (.A(reg_wdata[15]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_1 input22 (.A(reg_wdata[16]),
    .X(net22));
 sky130_fd_sc_hd__dlymetal6s2s_1 input23 (.A(reg_wdata[17]),
    .X(net23));
 sky130_fd_sc_hd__dlymetal6s2s_1 input24 (.A(reg_wdata[18]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(reg_wdata[19]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(reg_wdata[1]),
    .X(net26));
 sky130_fd_sc_hd__dlymetal6s2s_1 input27 (.A(reg_wdata[20]),
    .X(net27));
 sky130_fd_sc_hd__dlymetal6s2s_1 input28 (.A(reg_wdata[21]),
    .X(net28));
 sky130_fd_sc_hd__dlymetal6s2s_1 input29 (.A(reg_wdata[22]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(cfg_cska_usb[2]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input30 (.A(reg_wdata[23]),
    .X(net30));
 sky130_fd_sc_hd__dlymetal6s2s_1 input31 (.A(reg_wdata[28]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_1 input32 (.A(reg_wdata[29]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(reg_wdata[2]),
    .X(net33));
 sky130_fd_sc_hd__dlymetal6s2s_1 input34 (.A(reg_wdata[30]),
    .X(net34));
 sky130_fd_sc_hd__dlymetal6s2s_1 input35 (.A(reg_wdata[31]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_1 input36 (.A(reg_wdata[3]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(reg_wdata[4]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_1 input38 (.A(reg_wdata[5]),
    .X(net38));
 sky130_fd_sc_hd__dlymetal6s2s_1 input39 (.A(reg_wdata[6]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(cfg_cska_usb[3]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(reg_wdata[7]),
    .X(net40));
 sky130_fd_sc_hd__dlymetal6s2s_1 input41 (.A(reg_wdata[8]),
    .X(net41));
 sky130_fd_sc_hd__dlymetal6s2s_1 input42 (.A(reg_wdata[9]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(reg_wr),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(usb_in_dn),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(usb_in_dp),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 input46 (.A(usb_rstn),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(wbd_clk_int),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(reg_addr[0]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(reg_addr[1]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(reg_addr[2]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(reg_addr[3]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(reg_addr[4]),
    .X(net9));
 sky130_fd_sc_hd__buf_2 output48 (.A(net48),
    .X(reg_ack));
 sky130_fd_sc_hd__buf_2 output49 (.A(net49),
    .X(reg_rdata[0]));
 sky130_fd_sc_hd__buf_2 output50 (.A(net50),
    .X(reg_rdata[10]));
 sky130_fd_sc_hd__buf_2 output51 (.A(net51),
    .X(reg_rdata[11]));
 sky130_fd_sc_hd__buf_2 output52 (.A(net52),
    .X(reg_rdata[12]));
 sky130_fd_sc_hd__buf_2 output53 (.A(net53),
    .X(reg_rdata[13]));
 sky130_fd_sc_hd__buf_2 output54 (.A(net54),
    .X(reg_rdata[14]));
 sky130_fd_sc_hd__buf_2 output55 (.A(net55),
    .X(reg_rdata[15]));
 sky130_fd_sc_hd__buf_2 output56 (.A(net56),
    .X(reg_rdata[16]));
 sky130_fd_sc_hd__buf_2 output57 (.A(net57),
    .X(reg_rdata[17]));
 sky130_fd_sc_hd__buf_2 output58 (.A(net58),
    .X(reg_rdata[18]));
 sky130_fd_sc_hd__buf_2 output59 (.A(net59),
    .X(reg_rdata[19]));
 sky130_fd_sc_hd__buf_2 output60 (.A(net60),
    .X(reg_rdata[1]));
 sky130_fd_sc_hd__buf_2 output61 (.A(net61),
    .X(reg_rdata[20]));
 sky130_fd_sc_hd__buf_2 output62 (.A(net62),
    .X(reg_rdata[21]));
 sky130_fd_sc_hd__buf_2 output63 (.A(net63),
    .X(reg_rdata[22]));
 sky130_fd_sc_hd__buf_2 output64 (.A(net64),
    .X(reg_rdata[23]));
 sky130_fd_sc_hd__buf_2 output65 (.A(net65),
    .X(reg_rdata[24]));
 sky130_fd_sc_hd__buf_2 output66 (.A(net66),
    .X(reg_rdata[25]));
 sky130_fd_sc_hd__buf_2 output67 (.A(net67),
    .X(reg_rdata[26]));
 sky130_fd_sc_hd__buf_2 output68 (.A(net68),
    .X(reg_rdata[27]));
 sky130_fd_sc_hd__buf_2 output69 (.A(net69),
    .X(reg_rdata[28]));
 sky130_fd_sc_hd__buf_2 output70 (.A(net70),
    .X(reg_rdata[29]));
 sky130_fd_sc_hd__buf_2 output71 (.A(net71),
    .X(reg_rdata[2]));
 sky130_fd_sc_hd__buf_2 output72 (.A(net72),
    .X(reg_rdata[30]));
 sky130_fd_sc_hd__buf_2 output73 (.A(net73),
    .X(reg_rdata[31]));
 sky130_fd_sc_hd__buf_2 output74 (.A(net74),
    .X(reg_rdata[3]));
 sky130_fd_sc_hd__buf_2 output75 (.A(net75),
    .X(reg_rdata[4]));
 sky130_fd_sc_hd__buf_2 output76 (.A(net76),
    .X(reg_rdata[5]));
 sky130_fd_sc_hd__buf_2 output77 (.A(net77),
    .X(reg_rdata[6]));
 sky130_fd_sc_hd__buf_2 output78 (.A(net78),
    .X(reg_rdata[7]));
 sky130_fd_sc_hd__buf_2 output79 (.A(net79),
    .X(reg_rdata[8]));
 sky130_fd_sc_hd__buf_2 output80 (.A(net80),
    .X(reg_rdata[9]));
 sky130_fd_sc_hd__buf_2 output81 (.A(net81),
    .X(usb_intr_o));
 sky130_fd_sc_hd__buf_2 output82 (.A(net82),
    .X(usb_out_dn));
 sky130_fd_sc_hd__buf_2 output83 (.A(net83),
    .X(usb_out_dp));
 sky130_fd_sc_hd__buf_2 output84 (.A(net84),
    .X(usb_out_tx_oen));
 sky130_fd_sc_hd__buf_2 output85 (.A(net85),
    .X(wbd_clk_usb));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly0  (.A(\u_skew_usb.clk_inbuf ),
    .X(\u_skew_usb.clkbuf_1.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly1  (.A(\u_skew_usb.clkbuf_1.X1 ),
    .X(\u_skew_usb.clkbuf_1.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly2  (.A(\u_skew_usb.clkbuf_1.X2 ),
    .X(\u_skew_usb.clkbuf_1.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_1.u_dly3  (.A(\u_skew_usb.clkbuf_1.X3 ),
    .X(\u_skew_usb.clk_d1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly0  (.A(\u_skew_usb.clk_d9 ),
    .X(\u_skew_usb.clkbuf_10.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly1  (.A(\u_skew_usb.clkbuf_10.X1 ),
    .X(\u_skew_usb.clkbuf_10.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly2  (.A(\u_skew_usb.clkbuf_10.X2 ),
    .X(\u_skew_usb.clkbuf_10.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_10.u_dly3  (.A(\u_skew_usb.clkbuf_10.X3 ),
    .X(\u_skew_usb.clk_d10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly0  (.A(\u_skew_usb.clk_d10 ),
    .X(\u_skew_usb.clkbuf_11.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly1  (.A(\u_skew_usb.clkbuf_11.X1 ),
    .X(\u_skew_usb.clkbuf_11.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly2  (.A(\u_skew_usb.clkbuf_11.X2 ),
    .X(\u_skew_usb.clkbuf_11.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_11.u_dly3  (.A(\u_skew_usb.clkbuf_11.X3 ),
    .X(\u_skew_usb.clk_d11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly0  (.A(\u_skew_usb.clk_d11 ),
    .X(\u_skew_usb.clkbuf_12.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly1  (.A(\u_skew_usb.clkbuf_12.X1 ),
    .X(\u_skew_usb.clkbuf_12.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly2  (.A(\u_skew_usb.clkbuf_12.X2 ),
    .X(\u_skew_usb.clkbuf_12.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_12.u_dly3  (.A(\u_skew_usb.clkbuf_12.X3 ),
    .X(\u_skew_usb.clk_d12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly0  (.A(\u_skew_usb.clk_d12 ),
    .X(\u_skew_usb.clkbuf_13.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly1  (.A(\u_skew_usb.clkbuf_13.X1 ),
    .X(\u_skew_usb.clkbuf_13.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly2  (.A(\u_skew_usb.clkbuf_13.X2 ),
    .X(\u_skew_usb.clkbuf_13.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_13.u_dly3  (.A(\u_skew_usb.clkbuf_13.X3 ),
    .X(\u_skew_usb.clk_d13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly0  (.A(\u_skew_usb.clk_d13 ),
    .X(\u_skew_usb.clkbuf_14.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly1  (.A(\u_skew_usb.clkbuf_14.X1 ),
    .X(\u_skew_usb.clkbuf_14.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly2  (.A(\u_skew_usb.clkbuf_14.X2 ),
    .X(\u_skew_usb.clkbuf_14.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_14.u_dly3  (.A(\u_skew_usb.clkbuf_14.X3 ),
    .X(\u_skew_usb.clk_d14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly0  (.A(\u_skew_usb.clk_d14 ),
    .X(\u_skew_usb.clkbuf_15.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly1  (.A(\u_skew_usb.clkbuf_15.X1 ),
    .X(\u_skew_usb.clkbuf_15.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly2  (.A(\u_skew_usb.clkbuf_15.X2 ),
    .X(\u_skew_usb.clkbuf_15.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_15.u_dly3  (.A(\u_skew_usb.clkbuf_15.X3 ),
    .X(\u_skew_usb.clk_d15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly0  (.A(\u_skew_usb.clk_d1 ),
    .X(\u_skew_usb.clkbuf_2.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly1  (.A(\u_skew_usb.clkbuf_2.X1 ),
    .X(\u_skew_usb.clkbuf_2.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly2  (.A(\u_skew_usb.clkbuf_2.X2 ),
    .X(\u_skew_usb.clkbuf_2.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_2.u_dly3  (.A(\u_skew_usb.clkbuf_2.X3 ),
    .X(\u_skew_usb.clk_d2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly0  (.A(\u_skew_usb.clk_d2 ),
    .X(\u_skew_usb.clkbuf_3.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly1  (.A(\u_skew_usb.clkbuf_3.X1 ),
    .X(\u_skew_usb.clkbuf_3.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly2  (.A(\u_skew_usb.clkbuf_3.X2 ),
    .X(\u_skew_usb.clkbuf_3.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_3.u_dly3  (.A(\u_skew_usb.clkbuf_3.X3 ),
    .X(\u_skew_usb.clk_d3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly0  (.A(\u_skew_usb.clk_d3 ),
    .X(\u_skew_usb.clkbuf_4.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly1  (.A(\u_skew_usb.clkbuf_4.X1 ),
    .X(\u_skew_usb.clkbuf_4.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly2  (.A(\u_skew_usb.clkbuf_4.X2 ),
    .X(\u_skew_usb.clkbuf_4.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_4.u_dly3  (.A(\u_skew_usb.clkbuf_4.X3 ),
    .X(\u_skew_usb.clk_d4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly0  (.A(\u_skew_usb.clk_d4 ),
    .X(\u_skew_usb.clkbuf_5.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly1  (.A(\u_skew_usb.clkbuf_5.X1 ),
    .X(\u_skew_usb.clkbuf_5.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly2  (.A(\u_skew_usb.clkbuf_5.X2 ),
    .X(\u_skew_usb.clkbuf_5.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_5.u_dly3  (.A(\u_skew_usb.clkbuf_5.X3 ),
    .X(\u_skew_usb.clk_d5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly0  (.A(\u_skew_usb.clk_d5 ),
    .X(\u_skew_usb.clkbuf_6.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly1  (.A(\u_skew_usb.clkbuf_6.X1 ),
    .X(\u_skew_usb.clkbuf_6.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly2  (.A(\u_skew_usb.clkbuf_6.X2 ),
    .X(\u_skew_usb.clkbuf_6.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_6.u_dly3  (.A(\u_skew_usb.clkbuf_6.X3 ),
    .X(\u_skew_usb.clk_d6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly0  (.A(\u_skew_usb.clk_d6 ),
    .X(\u_skew_usb.clkbuf_7.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly1  (.A(\u_skew_usb.clkbuf_7.X1 ),
    .X(\u_skew_usb.clkbuf_7.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly2  (.A(\u_skew_usb.clkbuf_7.X2 ),
    .X(\u_skew_usb.clkbuf_7.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_7.u_dly3  (.A(\u_skew_usb.clkbuf_7.X3 ),
    .X(\u_skew_usb.clk_d7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly0  (.A(\u_skew_usb.clk_d7 ),
    .X(\u_skew_usb.clkbuf_8.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly1  (.A(\u_skew_usb.clkbuf_8.X1 ),
    .X(\u_skew_usb.clkbuf_8.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly2  (.A(\u_skew_usb.clkbuf_8.X2 ),
    .X(\u_skew_usb.clkbuf_8.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_8.u_dly3  (.A(\u_skew_usb.clkbuf_8.X3 ),
    .X(\u_skew_usb.clk_d8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly0  (.A(\u_skew_usb.clk_d8 ),
    .X(\u_skew_usb.clkbuf_9.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly1  (.A(\u_skew_usb.clkbuf_9.X1 ),
    .X(\u_skew_usb.clkbuf_9.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly2  (.A(\u_skew_usb.clkbuf_9.X2 ),
    .X(\u_skew_usb.clkbuf_9.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.clkbuf_9.u_dly3  (.A(\u_skew_usb.clkbuf_9.X3 ),
    .X(\u_skew_usb.clk_d9 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_clkbuf_in.u_buf  (.A(net47),
    .X(\u_skew_usb.clk_inbuf ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_clkbuf_out.u_buf  (.A(\u_skew_usb.d30 ),
    .X(net85));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_00.genblk1.u_mux  (.A0(\u_skew_usb.in0 ),
    .A1(\u_skew_usb.in1 ),
    .S(net1),
    .X(\u_skew_usb.d00 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_01.genblk1.u_mux  (.A0(\u_skew_usb.in2 ),
    .A1(\u_skew_usb.in3 ),
    .S(net1),
    .X(\u_skew_usb.d01 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_02.genblk1.u_mux  (.A0(\u_skew_usb.in4 ),
    .A1(\u_skew_usb.in5 ),
    .S(net1),
    .X(\u_skew_usb.d02 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_03.genblk1.u_mux  (.A0(\u_skew_usb.in6 ),
    .A1(\u_skew_usb.in7 ),
    .S(net1),
    .X(\u_skew_usb.d03 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_04.genblk1.u_mux  (.A0(\u_skew_usb.in8 ),
    .A1(\u_skew_usb.in9 ),
    .S(net1),
    .X(\u_skew_usb.d04 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_05.genblk1.u_mux  (.A0(\u_skew_usb.in10 ),
    .A1(\u_skew_usb.in11 ),
    .S(net1),
    .X(\u_skew_usb.d05 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_06.genblk1.u_mux  (.A0(\u_skew_usb.in12 ),
    .A1(\u_skew_usb.in13 ),
    .S(net1),
    .X(\u_skew_usb.d06 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_07.genblk1.u_mux  (.A0(\u_skew_usb.in14 ),
    .A1(\u_skew_usb.in15 ),
    .S(net1),
    .X(\u_skew_usb.d07 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_10.genblk1.u_mux  (.A0(\u_skew_usb.d00 ),
    .A1(\u_skew_usb.d01 ),
    .S(net2),
    .X(\u_skew_usb.d10 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_11.genblk1.u_mux  (.A0(\u_skew_usb.d02 ),
    .A1(\u_skew_usb.d03 ),
    .S(net2),
    .X(\u_skew_usb.d11 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_12.genblk1.u_mux  (.A0(\u_skew_usb.d04 ),
    .A1(\u_skew_usb.d05 ),
    .S(net2),
    .X(\u_skew_usb.d12 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_13.genblk1.u_mux  (.A0(\u_skew_usb.d06 ),
    .A1(\u_skew_usb.d07 ),
    .S(net2),
    .X(\u_skew_usb.d13 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_20.genblk1.u_mux  (.A0(\u_skew_usb.d10 ),
    .A1(\u_skew_usb.d11 ),
    .S(net3),
    .X(\u_skew_usb.d20 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_21.genblk1.u_mux  (.A0(\u_skew_usb.d12 ),
    .A1(\u_skew_usb.d13 ),
    .S(net3),
    .X(\u_skew_usb.d21 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_usb.u_mux_level_30.genblk1.u_mux  (.A0(\u_skew_usb.d20 ),
    .A1(\u_skew_usb.d21 ),
    .S(net4),
    .X(\u_skew_usb.d30 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_0.u_buf  (.A(\u_skew_usb.clk_inbuf ),
    .X(\u_skew_usb.in0 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_1.u_buf  (.A(\u_skew_usb.clk_d1 ),
    .X(\u_skew_usb.in1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_10.u_buf  (.A(\u_skew_usb.clk_d10 ),
    .X(\u_skew_usb.in10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_11.u_buf  (.A(\u_skew_usb.clk_d11 ),
    .X(\u_skew_usb.in11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_12.u_buf  (.A(\u_skew_usb.clk_d12 ),
    .X(\u_skew_usb.in12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_13.u_buf  (.A(\u_skew_usb.clk_d13 ),
    .X(\u_skew_usb.in13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_14.u_buf  (.A(\u_skew_usb.clk_d14 ),
    .X(\u_skew_usb.in14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_15.u_buf  (.A(\u_skew_usb.clk_d15 ),
    .X(\u_skew_usb.in15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_2.u_buf  (.A(\u_skew_usb.clk_d2 ),
    .X(\u_skew_usb.in2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_3.u_buf  (.A(\u_skew_usb.clk_d3 ),
    .X(\u_skew_usb.in3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_4.u_buf  (.A(\u_skew_usb.clk_d4 ),
    .X(\u_skew_usb.in4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_5.u_buf  (.A(\u_skew_usb.clk_d5 ),
    .X(\u_skew_usb.in5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_6.u_buf  (.A(\u_skew_usb.clk_d6 ),
    .X(\u_skew_usb.in6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_7.u_buf  (.A(\u_skew_usb.clk_d7 ),
    .X(\u_skew_usb.in7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_8.u_buf  (.A(\u_skew_usb.clk_d8 ),
    .X(\u_skew_usb.in8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_usb.u_tap_9.u_buf  (.A(\u_skew_usb.clk_d9 ),
    .X(\u_skew_usb.in9 ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._06_  (.A(\u_usb_host.u_async_wb.PendingRd ),
    .Y(\u_usb_host.u_async_wb._02_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._07_  (.A(\u_usb_host.u_async_wb.m_resp_rd_empty ),
    .Y(\u_usb_host.u_async_wb.m_resp_rd_en ));
 sky130_fd_sc_hd__or4b_2 \u_usb_host.u_async_wb._08_  (.A(\u_usb_host.u_async_wb.m_cmd_wr_full ),
    .B(\u_usb_host.u_async_wb.m_cmd_wr_afull ),
    .C(\u_usb_host.u_async_wb.PendingRd ),
    .D_N(\u_usb_host.u_async_wb.wbm_cyc_i ),
    .X(\u_usb_host.u_async_wb._03_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb._09_  (.A(\u_usb_host.u_async_wb._03_ ),
    .Y(\u_usb_host.u_async_wb.m_cmd_wr_en ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb._10_  (.A(net43),
    .B(\u_usb_host.u_async_wb._03_ ),
    .Y(\u_usb_host.u_async_wb._00_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_async_wb._11_  (.A(net43),
    .B(\u_usb_host.u_async_wb.m_resp_rd_empty ),
    .C_N(\u_usb_host.u_async_wb.wbm_cyc_i ),
    .X(\u_usb_host.u_async_wb._04_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_async_wb._12_  (.A1(net43),
    .A2(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .B1_N(\u_usb_host.u_async_wb._04_ ),
    .X(net48));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_async_wb._13_  (.A1(net43),
    .A2(\u_usb_host.u_async_wb._03_ ),
    .B1(\u_usb_host.u_async_wb._04_ ),
    .B2(\u_usb_host.u_async_wb._02_ ),
    .Y(\u_usb_host.u_async_wb._01_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._14_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[36] ),
    .X(\u_usb_host.reg_wr ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._19_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[4] ),
    .X(\u_usb_host.reg_wdata[0] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._20_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[5] ),
    .X(\u_usb_host.reg_wdata[1] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._21_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[6] ),
    .X(\u_usb_host.reg_wdata[2] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._22_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[7] ),
    .X(\u_usb_host.reg_wdata[3] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._23_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[8] ),
    .X(\u_usb_host.reg_wdata[4] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._24_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[9] ),
    .X(\u_usb_host.reg_wdata[5] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._25_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[10] ),
    .X(\u_usb_host.reg_wdata[6] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._26_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[11] ),
    .X(\u_usb_host.reg_wdata[7] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._27_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[12] ),
    .X(\u_usb_host.reg_wdata[8] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._28_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[13] ),
    .X(\u_usb_host.reg_wdata[9] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._29_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[14] ),
    .X(\u_usb_host.reg_wdata[10] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._30_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[15] ),
    .X(\u_usb_host.reg_wdata[11] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._31_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[16] ),
    .X(\u_usb_host.reg_wdata[12] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._32_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[17] ),
    .X(\u_usb_host.reg_wdata[13] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._33_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[18] ),
    .X(\u_usb_host.reg_wdata[14] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._34_  (.A_N(net110),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[19] ),
    .X(\u_usb_host.reg_wdata[15] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._35_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[20] ),
    .X(\u_usb_host.reg_wdata[16] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._36_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[21] ),
    .X(\u_usb_host.reg_wdata[17] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._37_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[22] ),
    .X(\u_usb_host.reg_wdata[18] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._38_  (.A_N(net109),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[23] ),
    .X(\u_usb_host.reg_wdata[19] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._39_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[24] ),
    .X(\u_usb_host.reg_wdata[20] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._40_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[25] ),
    .X(\u_usb_host.reg_wdata[21] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._41_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[26] ),
    .X(\u_usb_host.reg_wdata[22] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._42_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[27] ),
    .X(\u_usb_host.reg_wdata[23] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._47_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[32] ),
    .X(\u_usb_host.reg_wdata[28] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._48_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[33] ),
    .X(\u_usb_host.reg_wdata[29] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._49_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[34] ),
    .X(\u_usb_host.reg_wdata[30] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._50_  (.A_N(net108),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[35] ),
    .X(\u_usb_host.reg_wdata[31] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._51_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[37] ),
    .X(\u_usb_host.reg_addr[0] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._52_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[38] ),
    .X(\u_usb_host.reg_addr[1] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._53_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[39] ),
    .X(\u_usb_host.reg_addr[2] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._54_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[40] ),
    .X(\u_usb_host.reg_addr[3] ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_async_wb._55_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[41] ),
    .X(\u_usb_host.reg_addr[4] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_async_wb._56_  (.A_N(net107),
    .B(\u_usb_host.u_async_wb.s_cmd_rd_data[42] ),
    .X(\u_usb_host.reg_addr[5] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb._57_  (.A(net108),
    .B(\u_usb_host.u_async_wb.wbs_ack_f ),
    .Y(\u_usb_host.u_async_wb.wbs_cyc_o ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_async_wb._58_  (.A_N(\u_usb_host.u_async_wb.s_resp_wr_full ),
    .B_N(\u_usb_host.reg_wr ),
    .C(\u_usb_host.u_async_wb.wbs_cyc_o ),
    .D(\u_usb_host.reg_ack ),
    .X(\u_usb_host.u_async_wb.s_resp_wr_en ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb._59_  (.CLK(\u_usb_host.u_async_wb._05_ ),
    .D(\u_usb_host.u_async_wb._00_ ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.PendingRd ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb._60_  (.CLK(clknet_leaf_1_usb_clk),
    .D(\u_usb_host.reg_ack ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_async_wb.wbs_ack_f ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb._61_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb._01_ ),
    .GCLK(\u_usb_host.u_async_wb._05_ ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_async_wb._62_  (.A(\u_usb_host.u_async_wb.wbs_cyc_o ),
    .X(\u_usb_host.reg_cs ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._043_  (.A(net531),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._002_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_cmd_if._044_  (.A(net535),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._045_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._000_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_cmd_if._046_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_cmd_if._047_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._008_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_async_wb.u_cmd_if._048_  (.A(net531),
    .B(net535),
    .X(\u_usb_host.u_async_wb.u_cmd_if._009_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._049_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ),
    .B(net535),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._010_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_cmd_if._050_  (.A(\u_usb_host.u_async_wb.u_cmd_if._009_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._010_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._051_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_async_wb.u_cmd_if._052_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._011_ ));
 sky130_fd_sc_hd__xnor2_2 \u_usb_host.u_async_wb.u_cmd_if._053_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._011_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._012_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_async_wb.u_cmd_if._054_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._013_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._055_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._011_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._014_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_async_wb.u_cmd_if._056_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._014_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._015_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._057_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._016_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._058_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._017_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._059_  (.A(\u_usb_host.u_async_wb.u_cmd_if._015_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._016_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._017_ ),
    .X(\u_usb_host.u_async_wb.m_cmd_wr_full ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_async_wb.u_cmd_if._060_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .C_N(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._018_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._061_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._019_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._062_  (.A1(\u_usb_host.u_async_wb.u_cmd_if._013_ ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._018_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._016_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._020_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._063_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._012_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._014_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._021_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_async_wb.u_cmd_if._064_  (.A1(\u_usb_host.u_async_wb.u_cmd_if._013_ ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if._016_ ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if._018_ ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._021_ ),
    .C1(\u_usb_host.u_async_wb.u_cmd_if._015_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._022_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_cmd_if._065_  (.A(\u_usb_host.u_async_wb.u_cmd_if._020_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._022_ ),
    .Y(\u_usb_host.u_async_wb.m_cmd_wr_afull ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_cmd_if._066_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._023_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._067_  (.A(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._023_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._024_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_async_wb.u_cmd_if._068_  (.A(net535),
    .B(\u_usb_host.u_async_wb.u_cmd_if._024_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._025_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_async_wb.u_cmd_if._069_  (.A(net539),
    .B(\u_usb_host.u_async_wb.u_cmd_if._024_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._026_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._070_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._023_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._027_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_cmd_if._073_  (.A0(\u_usb_host.u_async_wb.u_cmd_if._008_ ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ),
    .S(\u_usb_host.u_async_wb.u_cmd_if._002_ ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._030_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._074_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._030_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._031_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_async_wb.u_cmd_if._076_  (.A(\u_usb_host.u_async_wb.u_cmd_if._025_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._026_ ),
    .C(\u_usb_host.u_async_wb.u_cmd_if._027_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._031_ ),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_empty ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._078_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._019_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_cmd_if._079_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._033_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._080_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._033_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._001_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_cmd_if._081_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if._010_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_cmd_if._082_  (.A(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._034_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_async_wb.u_cmd_if._083_  (.A1(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .B1(\u_usb_host.u_async_wb.u_cmd_if._034_ ),
    .Y(\u_usb_host.u_async_wb.u_cmd_if._003_ ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._088_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[4] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._089_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ),
    .S0(net538),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[5] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._090_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ),
    .S0(net538),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[6] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._091_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ),
    .S0(net536),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[7] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._092_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[8] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._093_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[9] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._094_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ),
    .S0(net537),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[10] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._095_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ),
    .S0(net538),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[11] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._096_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ),
    .S0(net538),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[12] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._097_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[13] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._098_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ),
    .S0(net538),
    .S1(net534),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[14] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._099_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[15] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._100_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[16] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._101_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ),
    .S0(net538),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[17] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._102_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ),
    .S0(net538),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[18] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._103_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[19] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._104_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[20] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._105_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[21] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._106_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[22] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._107_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[23] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._108_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[24] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._109_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[25] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._110_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ),
    .S0(net539),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[26] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._111_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[27] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._116_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ),
    .S0(net539),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[32] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._117_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[33] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._118_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ),
    .S0(net537),
    .S1(net533),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[34] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._119_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[35] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._120_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[36] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._121_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[37] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._122_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[38] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._123_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[39] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._124_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[40] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._125_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ),
    .S0(net535),
    .S1(net531),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[41] ));
 sky130_fd_sc_hd__mux4_1 \u_usb_host.u_async_wb.u_cmd_if._126_  (.A0(\u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ),
    .A1(\u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ),
    .A2(\u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ),
    .A3(\u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ),
    .S0(net536),
    .S1(net532),
    .X(\u_usb_host.u_async_wb.s_cmd_rd_data[42] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._127_  (.A(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._006_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._128_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._005_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._129_  (.A(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._004_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_async_wb.u_cmd_if._130_  (.A(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .B(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .C(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .X(\u_usb_host.u_async_wb.u_cmd_if._007_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._135_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._136_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._137_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._138_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._139_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._140_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._141_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._142_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._143_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._144_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._145_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._146_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._147_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._148_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._149_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._150_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._151_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._152_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._153_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._154_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._155_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._156_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._157_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._158_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._163_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._164_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._165_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._166_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._167_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._168_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._169_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._170_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._171_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._172_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._173_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._041_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[1][42] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._178_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._179_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._180_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._181_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._182_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._183_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._184_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._185_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._186_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._187_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._188_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._189_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._190_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._191_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._192_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._193_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._194_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._195_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._196_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._197_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._198_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._199_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._200_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._201_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._206_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._207_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._208_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._209_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._210_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._211_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._212_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._213_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._214_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._215_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._216_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._040_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[2][42] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._221_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._222_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._223_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._224_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._225_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._226_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._227_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._228_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._229_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._230_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._231_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._232_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._233_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._234_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._235_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._236_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._237_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._238_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._239_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._240_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._241_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._242_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._243_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._244_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._249_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._250_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._251_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._252_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._253_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._254_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._255_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._256_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._257_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._258_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._259_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._039_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[3][42] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._260_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._002_ ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._261_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._003_ ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._262_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._038_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._267_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net15),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._268_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net26),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._269_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net33),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._270_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net36),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._271_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net37),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._272_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net38),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._273_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net39),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._274_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net40),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._275_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net41),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._276_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net42),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._277_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net16),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._278_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net17),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._279_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net18),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._280_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net19),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._281_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net20),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._282_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net21),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._283_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net22),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._284_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net23),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._285_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net24),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._286_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net25),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._287_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net27),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._288_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net28),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._289_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net29),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._290_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net30),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._295_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net31),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][32] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._296_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net32),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][33] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._297_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net34),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][34] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._298_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net35),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][35] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._299_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net43),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][36] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._300_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net5),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][37] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._301_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net6),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][38] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._302_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net7),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][39] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._303_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net8),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][40] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._304_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net9),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][41] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_cmd_if._305_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_cmd_if._042_ ),
    .D(net10),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.mem[0][42] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_async_wb.u_cmd_if._306_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[0] ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_cmd_if._307_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[1] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._308_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._036_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._309_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._000_ ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._310_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if._001_ ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._311_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._037_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.wr_ptr_inc[2] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._312_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[0] ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_cmd_if._313_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[1] ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._314_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_cmd_if._035_ ),
    .D(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr_inc[2] ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._315_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[0] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._316_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[1] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._317_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_rd_ptr[2] ),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._318_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net674),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._319_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net673),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._320_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net658),
    .RESET_B(net365),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._321_  (.CLK(clknet_leaf_59_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[0] ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._322_  (.CLK(clknet_leaf_59_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[1] ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._323_  (.CLK(clknet_leaf_59_usb_clk),
    .D(\u_usb_host.u_async_wb.u_cmd_if.grey_wr_ptr[2] ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._324_  (.CLK(clknet_leaf_59_usb_clk),
    .D(net655),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._325_  (.CLK(clknet_leaf_59_usb_clk),
    .D(net657),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_cmd_if._326_  (.CLK(clknet_leaf_59_usb_clk),
    .D(net656),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_cmd_if.sync_wr_ptr[2] ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._327_  (.CLK(clknet_leaf_2_usb_clk),
    .GATE(\u_usb_host.reg_ack ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._035_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._328_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._036_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._329_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_cmd_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._037_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_cmd_if._330_  (.CLK(clknet_leaf_2_usb_clk),
    .GATE(\u_usb_host.reg_ack ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._038_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._331_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._004_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._039_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._332_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._005_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._040_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._333_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._006_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._041_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_cmd_if._334_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.u_cmd_if._007_ ),
    .GCLK(\u_usb_host.u_async_wb.u_cmd_if._042_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_resp_if._020_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._012_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_resp_if._021_  (.A(net530),
    .Y(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_async_wb.u_resp_if._022_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_async_wb.u_resp_if._023_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._010_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._024_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._025_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(net530),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._026_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._002_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._027_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if._002_ ),
    .X(\u_usb_host.u_async_wb.u_resp_if._003_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._028_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if._004_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_resp_if._029_  (.A1(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .A2(\u_usb_host.u_async_wb.u_resp_if._002_ ),
    .B1(\u_usb_host.u_async_wb.u_resp_if._004_ ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._005_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_resp_if._030_  (.A(\u_usb_host.u_async_wb.u_resp_if._003_ ),
    .B(\u_usb_host.u_async_wb.u_resp_if._005_ ),
    .Y(\u_usb_host.u_async_wb.s_resp_wr_full ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._032_  (.A(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._006_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._033_  (.A(net530),
    .B(\u_usb_host.u_async_wb.u_resp_if._006_ ),
    .X(\u_usb_host.u_async_wb.u_resp_if._007_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_async_wb.u_resp_if._034_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._008_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_async_wb.u_resp_if._035_  (.A1(net530),
    .A2(\u_usb_host.u_async_wb.u_resp_if._006_ ),
    .B1(\u_usb_host.u_async_wb.u_resp_if._008_ ),
    .Y(\u_usb_host.u_async_wb.u_resp_if._009_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_async_wb.u_resp_if._036_  (.A(\u_usb_host.u_async_wb.u_resp_if._007_ ),
    .B(\u_usb_host.u_async_wb.u_resp_if._009_ ),
    .Y(\u_usb_host.u_async_wb.m_resp_rd_empty ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._038_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][0] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][0] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._039_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][1] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][1] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[1] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._040_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][2] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][2] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[2] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._041_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][3] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][3] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[3] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._042_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][4] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][4] ),
    .S(net569),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[4] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._043_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][5] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][5] ),
    .S(net569),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[5] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._044_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][6] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][6] ),
    .S(net569),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[6] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._045_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][7] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][7] ),
    .S(net569),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[7] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._046_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][8] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][8] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[8] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._047_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][9] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][9] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[9] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._048_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][10] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][10] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[10] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._049_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][11] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][11] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[11] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._050_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][12] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][12] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[12] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._051_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][13] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][13] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[13] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._052_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][14] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][14] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[14] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._053_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][15] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][15] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[15] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._054_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][16] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][16] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[16] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._055_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][17] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][17] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[17] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._056_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][18] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][18] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[18] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._057_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][19] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][19] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[19] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._058_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][20] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][20] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[20] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._059_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][21] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][21] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[21] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._060_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][22] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][22] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[22] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._061_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][23] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][23] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[23] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._062_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][24] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][24] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[24] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._063_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][25] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][25] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[25] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._064_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][26] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][26] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[26] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._065_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][27] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][27] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[27] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._066_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][28] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][28] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[28] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._067_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][29] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][29] ),
    .S(net528),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[29] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._068_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][30] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][30] ),
    .S(net527),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[30] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_async_wb.u_resp_if._069_  (.A0(\u_usb_host.u_async_wb.u_resp_if.mem[0][31] ),
    .A1(\u_usb_host.u_async_wb.u_resp_if.mem[1][31] ),
    .S(net526),
    .X(\u_usb_host.u_async_wb.u_resp_if.rd_data[31] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._071_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .X(\u_usb_host.u_async_wb.u_resp_if._000_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_async_wb.u_resp_if._072_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ),
    .B(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .X(\u_usb_host.u_async_wb.u_resp_if._001_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._073_  (.A(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ),
    .B(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ),
    .X(\u_usb_host.u_async_wb.u_resp_if._011_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_async_wb.u_resp_if._074_  (.A(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ),
    .B(net530),
    .X(\u_usb_host.u_async_wb.u_resp_if._013_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._075_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net608),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._076_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net605),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._077_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net609),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._078_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net618),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._079_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net623),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._080_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net617),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._081_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net607),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._082_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net619),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._083_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net596),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._084_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net604),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._085_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net626),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._086_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net599),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._087_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net606),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._088_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net603),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._089_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net627),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._090_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net629),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._091_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net598),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._092_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net645),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._093_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net625),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._094_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net630),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._095_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net628),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._096_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net597),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._097_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net602),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._098_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net644),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._099_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net646),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._100_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net668),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._101_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net643),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._102_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net632),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._103_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net600),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][28] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._104_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net613),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][29] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._105_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net640),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][30] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._106_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._018_ ),
    .D(net610),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[1][31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._108_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[0] ),
    .RESET_B(net571),
    .Q(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._109_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._014_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.rd_ptr_inc[1] ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.rd_ptr[1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._110_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net608),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._111_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net605),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._112_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net609),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._113_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net618),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._114_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net623),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._115_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net617),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._116_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net607),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._117_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net619),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._118_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net596),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._119_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net604),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._120_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net626),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._121_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net599),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._122_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net606),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._123_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net603),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._124_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net627),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._125_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net629),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._126_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net598),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._127_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net645),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._128_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net625),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._129_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net630),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._130_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net628),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._131_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net597),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._132_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net602),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._133_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net644),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][23] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._134_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net646),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][24] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._135_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net668),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][25] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._136_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net643),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][26] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._137_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net632),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][27] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._138_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net600),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][28] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._139_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net613),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][29] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._140_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net640),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][30] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_async_wb.u_resp_if._141_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_async_wb.u_resp_if._019_ ),
    .D(net610),
    .Q(\u_usb_host.u_async_wb.u_resp_if.mem[0][31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._143_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._010_ ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._144_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._016_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._011_ ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._145_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._012_ ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._146_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._017_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if._013_ ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._147_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[0] ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_async_wb.u_resp_if._148_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_async_wb.u_resp_if._015_ ),
    .D(\u_usb_host.u_async_wb.u_resp_if.wr_ptr_inc[1] ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_async_wb.u_resp_if.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._149_  (.CLK(clknet_leaf_1_usb_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[0] ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._150_  (.CLK(clknet_leaf_1_usb_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_rd_ptr[1] ),
    .RESET_B(net368),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._151_  (.CLK(clknet_leaf_1_usb_clk),
    .D(net681),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._152_  (.CLK(clknet_leaf_1_usb_clk),
    .D(net679),
    .RESET_B(net367),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_rd_ptr_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._153_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[0] ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._154_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(\u_usb_host.u_async_wb.u_resp_if.grey_wr_ptr[1] ),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._155_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(net677),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_async_wb.u_resp_if._156_  (.CLK(clknet_1_1__leaf_app_clk),
    .D(net680),
    .RESET_B(net364),
    .Q(\u_usb_host.u_async_wb.u_resp_if.sync_wr_ptr_1[1] ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._157_  (.CLK(clknet_1_0__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_resp_rd_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._014_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._158_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._015_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._159_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_async_wb.s_resp_wr_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._016_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_async_wb.u_resp_if._160_  (.CLK(clknet_1_1__leaf_app_clk),
    .GATE(\u_usb_host.u_async_wb.m_resp_rd_en ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._017_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_resp_if._161_  (.CLK(clknet_leaf_7_usb_clk),
    .GATE(\u_usb_host.u_async_wb.u_resp_if._000_ ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._018_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_async_wb.u_resp_if._162_  (.CLK(clknet_leaf_7_usb_clk),
    .GATE(\u_usb_host.u_async_wb.u_resp_if._001_ ),
    .GCLK(\u_usb_host.u_async_wb.u_resp_if._019_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._203_  (.A(\u_usb_host.u_core.sof_time_q[0] ),
    .Y(\u_usb_host.u_core._007_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._204_  (.A(\u_usb_host.u_core.sof_time_q[12] ),
    .Y(\u_usb_host.u_core._061_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._205_  (.A(\u_usb_host.u_core.sof_time_q[14] ),
    .Y(\u_usb_host.u_core._062_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._206_  (.A(\u_usb_host.u_core.sof_value_q[0] ),
    .Y(\u_usb_host.u_core._050_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._207_  (.A(net614),
    .Y(\u_usb_host.u_core._026_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._208_  (.A(net682),
    .Y(\u_usb_host.u_core._002_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._209_  (.A(\u_usb_host.reg_addr[2] ),
    .Y(\u_usb_host.u_core._063_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core._210_  (.A(\u_usb_host.u_core.transfer_ack_w ),
    .Y(\u_usb_host.u_core._064_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._211_  (.A(\u_usb_host.u_core.sof_time_q[1] ),
    .B(\u_usb_host.u_core.sof_time_q[0] ),
    .C(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._065_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core._212_  (.A(\u_usb_host.u_core.sof_time_q[1] ),
    .B(\u_usb_host.u_core.sof_time_q[0] ),
    .C(\u_usb_host.u_core.sof_time_q[3] ),
    .D(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._066_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._213_  (.A(\u_usb_host.u_core.sof_time_q[14] ),
    .B(\u_usb_host.u_core.sof_time_q[15] ),
    .Y(\u_usb_host.u_core._067_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core._214_  (.A_N(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core.sof_time_q[14] ),
    .D(\u_usb_host.u_core.sof_time_q[15] ),
    .X(\u_usb_host.u_core._068_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core._215_  (.A_N(\u_usb_host.u_core.sof_time_q[8] ),
    .B_N(\u_usb_host.u_core.sof_time_q[12] ),
    .C(\u_usb_host.u_core.sof_time_q[13] ),
    .D(\u_usb_host.u_core.sof_time_q[9] ),
    .X(\u_usb_host.u_core._069_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core._216_  (.A_N(\u_usb_host.u_core.sof_time_q[5] ),
    .B_N(\u_usb_host.u_core.sof_time_q[7] ),
    .C(\u_usb_host.u_core.sof_time_q[6] ),
    .D(\u_usb_host.u_core.sof_time_q[4] ),
    .X(\u_usb_host.u_core._070_ ));
 sky130_fd_sc_hd__nand4_1 \u_usb_host.u_core._217_  (.A(\u_usb_host.u_core._066_ ),
    .B(\u_usb_host.u_core._068_ ),
    .C(\u_usb_host.u_core._069_ ),
    .D(\u_usb_host.u_core._070_ ),
    .Y(\u_usb_host.u_core._071_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._218_  (.A(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .B(net113),
    .Y(\u_usb_host.u_core._072_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core._219_  (.A(\u_usb_host.u_core._071_ ),
    .B(\u_usb_host.u_core._072_ ),
    .X(\u_usb_host.u_core._073_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._220_  (.A(\u_usb_host.u_core._073_ ),
    .Y(\u_usb_host.u_core.send_sof_w ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._221_  (.A(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .B(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .X(\u_usb_host.u_core._000_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._222_  (.A(\u_usb_host.u_core.usb_irq_ack_device_detect_out_w ),
    .B(\u_usb_host.u_core._000_ ),
    .X(\u_usb_host.u_core._045_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._223_  (.A(\u_usb_host.u_core.status_timeout_w ),
    .B(\u_usb_host.u_core.status_crc_err_w ),
    .X(\u_usb_host.u_core._001_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._224_  (.A_N(\u_usb_host.u_core.err_cond_q ),
    .B(\u_usb_host.u_core._001_ ),
    .X(\u_usb_host.u_core._004_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._225_  (.A(\u_usb_host.u_core.usb_irq_ack_err_out_w ),
    .B(\u_usb_host.u_core._004_ ),
    .X(\u_usb_host.u_core._044_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._226_  (.A(\u_usb_host.u_core.sof_irq_q ),
    .B(\u_usb_host.u_core.usb_irq_ack_sof_out_w ),
    .X(\u_usb_host.u_core._043_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._227_  (.A(\u_usb_host.u_core.status_tx_done_w ),
    .B(\u_usb_host.u_core.status_rx_done_w ),
    .X(\u_usb_host.u_core._003_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._228_  (.A(\u_usb_host.u_core.usb_irq_ack_done_out_w ),
    .B(\u_usb_host.u_core._003_ ),
    .X(\u_usb_host.u_core._042_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._229_  (.A(\u_usb_host.u_core.usb_ctrl_wr_q ),
    .B(\u_usb_host.u_core.utmi_rxerror_i ),
    .X(\u_usb_host.u_core._041_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_core._230_  (.A_N(\u_usb_host.u_core._071_ ),
    .B(\u_usb_host.u_core._072_ ),
    .Y(\u_usb_host.u_core._040_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core._231_  (.A1(\u_usb_host.u_core.sof_time_q[1] ),
    .A2(\u_usb_host.u_core.sof_time_q[0] ),
    .B1(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._074_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_core._232_  (.A1(\u_usb_host.u_core.sof_time_q[3] ),
    .A2(\u_usb_host.u_core.sof_time_q[4] ),
    .A3(\u_usb_host.u_core._074_ ),
    .B1(\u_usb_host.u_core.sof_time_q[6] ),
    .C1(\u_usb_host.u_core.sof_time_q[5] ),
    .X(\u_usb_host.u_core._075_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core._233_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core.sof_time_q[8] ),
    .C(\u_usb_host.u_core.sof_time_q[9] ),
    .D(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._076_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core._234_  (.A(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core.sof_time_q[14] ),
    .C(\u_usb_host.u_core.sof_time_q[15] ),
    .D(\u_usb_host.u_core._076_ ),
    .X(\u_usb_host.u_core._077_ ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_core._235_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core._075_ ),
    .D(\u_usb_host.u_core._077_ ),
    .Y(\u_usb_host.u_core._078_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._236_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._079_ ));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_core._237_  (.A1(\u_usb_host.u_core.sof_time_q[13] ),
    .A2(\u_usb_host.u_core._079_ ),
    .B1_N(\u_usb_host.u_core._067_ ),
    .X(\u_usb_host.u_core._080_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core._238_  (.A(\u_usb_host.u_core.sof_time_q[1] ),
    .B(\u_usb_host.u_core.sof_time_q[0] ),
    .C(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._081_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_core._239_  (.A1(\u_usb_host.u_core.sof_time_q[3] ),
    .A2(\u_usb_host.u_core.sof_time_q[5] ),
    .A3(\u_usb_host.u_core.sof_time_q[4] ),
    .A4(\u_usb_host.u_core._081_ ),
    .B1(\u_usb_host.u_core.sof_time_q[6] ),
    .X(\u_usb_host.u_core._082_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core._240_  (.A_N(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core.sof_time_q[9] ),
    .C(\u_usb_host.u_core.sof_time_q[8] ),
    .D(\u_usb_host.u_core.sof_time_q[7] ),
    .X(\u_usb_host.u_core._083_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._241_  (.A(\u_usb_host.u_core.sof_time_q[12] ),
    .B(\u_usb_host.u_core._068_ ),
    .C(\u_usb_host.u_core._082_ ),
    .D(\u_usb_host.u_core._083_ ),
    .X(\u_usb_host.u_core._084_ ));
 sky130_fd_sc_hd__o31ai_2 \u_usb_host.u_core._242_  (.A1(\u_usb_host.u_core._078_ ),
    .A2(\u_usb_host.u_core._080_ ),
    .A3(\u_usb_host.u_core._084_ ),
    .B1(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .Y(\u_usb_host.u_core._085_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._243_  (.A1(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .A2(net113),
    .A3(\u_usb_host.u_core._085_ ),
    .B1(\u_usb_host.u_core.send_sof_w ),
    .X(\u_usb_host.u_core._086_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._244_  (.A(\u_usb_host.u_core._002_ ),
    .B(\u_usb_host.u_core._086_ ),
    .X(\u_usb_host.u_core._039_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._245_  (.A1(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ),
    .A2(net113),
    .A3(\u_usb_host.u_core._085_ ),
    .B1(\u_usb_host.u_core.transfer_start_q ),
    .X(\u_usb_host.u_core._038_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core._246_  (.A_N(\u_usb_host.reg_addr[5] ),
    .B(\u_usb_host.reg_addr[4] ),
    .Y(\u_usb_host.u_core._087_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._247_  (.A(\u_usb_host.reg_addr[1] ),
    .B(\u_usb_host.reg_addr[0] ),
    .Y(\u_usb_host.u_core._088_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._248_  (.A(\u_usb_host.reg_addr[3] ),
    .B(\u_usb_host.u_core._088_ ),
    .Y(\u_usb_host.u_core._089_ ));
 sky130_fd_sc_hd__or3b_2 \u_usb_host.u_core._249_  (.A(\u_usb_host.u_core._089_ ),
    .B(\u_usb_host.reg_addr[2] ),
    .C_N(\u_usb_host.u_core.cfg_wr ),
    .X(\u_usb_host.u_core._090_ ));
 sky130_fd_sc_hd__nor2_4 \u_usb_host.u_core._250_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._090_ ),
    .Y(\u_usb_host.u_core._037_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core._251_  (.A(\u_usb_host.reg_addr[2] ),
    .B(\u_usb_host.u_core._087_ ),
    .C(\u_usb_host.u_core._089_ ),
    .Y(\u_usb_host.u_core._091_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._252_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core._037_ ),
    .X(\u_usb_host.u_core._036_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._253_  (.A_N(\u_usb_host.reg_ack ),
    .B(\u_usb_host.reg_cs ),
    .X(\u_usb_host.u_core._006_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._254_  (.A(\u_usb_host.reg_wr ),
    .B(\u_usb_host.u_core._006_ ),
    .X(\u_usb_host.u_core._047_ ));
 sky130_fd_sc_hd__or4_4 \u_usb_host.u_core._255_  (.A(\u_usb_host.reg_addr[1] ),
    .B(\u_usb_host.reg_addr[0] ),
    .C(\u_usb_host.reg_addr[2] ),
    .D(\u_usb_host.reg_addr[3] ),
    .X(\u_usb_host.u_core._092_ ));
 sky130_fd_sc_hd__or2_4 \u_usb_host.u_core._256_  (.A(\u_usb_host.reg_addr[5] ),
    .B(\u_usb_host.reg_addr[4] ),
    .X(\u_usb_host.u_core._093_ ));
 sky130_fd_sc_hd__nor2_8 \u_usb_host.u_core._257_  (.A(\u_usb_host.u_core._092_ ),
    .B(\u_usb_host.u_core._093_ ),
    .Y(\u_usb_host.u_core._094_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core._258_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._094_ ),
    .X(\u_usb_host.u_core._025_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core._259_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._092_ ),
    .Y(\u_usb_host.u_core._095_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._260_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._095_ ),
    .X(\u_usb_host.u_core._034_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_core._261_  (.A(\u_usb_host.u_core._063_ ),
    .B(\u_usb_host.reg_addr[3] ),
    .C_N(\u_usb_host.u_core._088_ ),
    .X(\u_usb_host.u_core._096_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._262_  (.A(\u_usb_host.u_core._087_ ),
    .B(\u_usb_host.u_core._096_ ),
    .Y(\u_usb_host.u_core._097_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._263_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(net92),
    .X(\u_usb_host.u_core._035_ ));
 sky130_fd_sc_hd__nor3b_4 \u_usb_host.u_core._264_  (.A(\u_usb_host.reg_addr[4] ),
    .B(\u_usb_host.u_core._092_ ),
    .C_N(\u_usb_host.reg_addr[5] ),
    .Y(\u_usb_host.u_core._098_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._265_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.u_core._098_ ),
    .X(\u_usb_host.u_core._031_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._266_  (.A(\u_usb_host.u_core._093_ ),
    .B(\u_usb_host.u_core._096_ ),
    .Y(\u_usb_host.u_core._099_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._267_  (.A(\u_usb_host.u_core.sof_time_q[8] ),
    .B(net89),
    .X(\u_usb_host.u_core.reg_rdata_r[24] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._268_  (.A(\u_usb_host.u_core.sof_time_q[9] ),
    .B(net89),
    .X(\u_usb_host.u_core.reg_rdata_r[25] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._269_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(net89),
    .X(\u_usb_host.u_core.reg_rdata_r[26] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._270_  (.A(\u_usb_host.u_core.sof_time_q[11] ),
    .B(net89),
    .X(\u_usb_host.u_core.reg_rdata_r[27] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._271_  (.A(\u_usb_host.u_core.sof_time_q[1] ),
    .B(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._014_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._272_  (.A1(\u_usb_host.u_core.sof_time_q[1] ),
    .A2(\u_usb_host.u_core.sof_time_q[0] ),
    .B1(\u_usb_host.u_core.sof_time_q[2] ),
    .Y(\u_usb_host.u_core._100_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._273_  (.A(\u_usb_host.u_core._065_ ),
    .B(\u_usb_host.u_core._100_ ),
    .Y(\u_usb_host.u_core._015_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._274_  (.A(\u_usb_host.u_core.sof_time_q[3] ),
    .B(\u_usb_host.u_core._065_ ),
    .Y(\u_usb_host.u_core._101_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._275_  (.A(\u_usb_host.u_core._066_ ),
    .B(\u_usb_host.u_core._101_ ),
    .Y(\u_usb_host.u_core._016_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._276_  (.A(\u_usb_host.u_core.sof_time_q[4] ),
    .B(\u_usb_host.u_core._066_ ),
    .X(\u_usb_host.u_core._017_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._277_  (.A(\u_usb_host.u_core.sof_time_q[5] ),
    .B(\u_usb_host.u_core.sof_time_q[4] ),
    .C(\u_usb_host.u_core._066_ ),
    .X(\u_usb_host.u_core._102_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._278_  (.A1(\u_usb_host.u_core.sof_time_q[4] ),
    .A2(\u_usb_host.u_core._066_ ),
    .B1(\u_usb_host.u_core.sof_time_q[5] ),
    .Y(\u_usb_host.u_core._103_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core._279_  (.A(\u_usb_host.u_core.send_sof_w ),
    .B(\u_usb_host.u_core._102_ ),
    .C(\u_usb_host.u_core._103_ ),
    .Y(\u_usb_host.u_core._018_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._280_  (.A(\u_usb_host.u_core.sof_time_q[5] ),
    .B(\u_usb_host.u_core.sof_time_q[4] ),
    .C(\u_usb_host.u_core.sof_time_q[6] ),
    .D(\u_usb_host.u_core._066_ ),
    .X(\u_usb_host.u_core._104_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._281_  (.A(\u_usb_host.u_core.send_sof_w ),
    .B(\u_usb_host.u_core._104_ ),
    .Y(\u_usb_host.u_core._105_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core._282_  (.A1(\u_usb_host.u_core.sof_time_q[6] ),
    .A2(\u_usb_host.u_core._102_ ),
    .B1(\u_usb_host.u_core._105_ ),
    .X(\u_usb_host.u_core._019_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._283_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core._104_ ),
    .Y(\u_usb_host.u_core._106_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._284_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core._104_ ),
    .X(\u_usb_host.u_core._107_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._285_  (.A(\u_usb_host.u_core._106_ ),
    .B(\u_usb_host.u_core._107_ ),
    .X(\u_usb_host.u_core._020_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core._286_  (.A(\u_usb_host.u_core.sof_time_q[8] ),
    .B(\u_usb_host.u_core._106_ ),
    .Y(\u_usb_host.u_core._021_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core._287_  (.A1(\u_usb_host.u_core.sof_time_q[7] ),
    .A2(\u_usb_host.u_core.sof_time_q[8] ),
    .A3(\u_usb_host.u_core._104_ ),
    .B1(\u_usb_host.u_core.sof_time_q[9] ),
    .X(\u_usb_host.u_core._108_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core._288_  (.A(\u_usb_host.u_core.sof_time_q[7] ),
    .B(\u_usb_host.u_core.sof_time_q[8] ),
    .C(\u_usb_host.u_core.sof_time_q[9] ),
    .D(\u_usb_host.u_core._104_ ),
    .X(\u_usb_host.u_core._109_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._289_  (.A(\u_usb_host.u_core._109_ ),
    .Y(\u_usb_host.u_core._110_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._290_  (.A(\u_usb_host.u_core._073_ ),
    .B(\u_usb_host.u_core._108_ ),
    .C(\u_usb_host.u_core._110_ ),
    .X(\u_usb_host.u_core._022_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._291_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core._109_ ),
    .X(\u_usb_host.u_core._008_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._292_  (.A1(\u_usb_host.u_core.sof_time_q[10] ),
    .A2(\u_usb_host.u_core._109_ ),
    .B1(\u_usb_host.u_core.sof_time_q[11] ),
    .X(\u_usb_host.u_core._111_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core._293_  (.A(\u_usb_host.u_core.sof_time_q[10] ),
    .B(\u_usb_host.u_core.sof_time_q[11] ),
    .C(\u_usb_host.u_core._109_ ),
    .Y(\u_usb_host.u_core._112_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._294_  (.A(\u_usb_host.u_core._073_ ),
    .B(\u_usb_host.u_core._111_ ),
    .C(\u_usb_host.u_core._112_ ),
    .X(\u_usb_host.u_core._009_ ));
 sky130_fd_sc_hd__a22oi_1 \u_usb_host.u_core._295_  (.A1(\u_usb_host.u_core._079_ ),
    .A2(\u_usb_host.u_core._109_ ),
    .B1(\u_usb_host.u_core._112_ ),
    .B2(\u_usb_host.u_core._061_ ),
    .Y(\u_usb_host.u_core._010_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._296_  (.A1(\u_usb_host.u_core._079_ ),
    .A2(\u_usb_host.u_core._109_ ),
    .B1(\u_usb_host.u_core.sof_time_q[13] ),
    .X(\u_usb_host.u_core._113_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core._297_  (.A(\u_usb_host.u_core.sof_time_q[13] ),
    .B(\u_usb_host.u_core._079_ ),
    .C(\u_usb_host.u_core._109_ ),
    .Y(\u_usb_host.u_core._114_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._298_  (.A(\u_usb_host.u_core._073_ ),
    .B(\u_usb_host.u_core._113_ ),
    .C(\u_usb_host.u_core._114_ ),
    .X(\u_usb_host.u_core._011_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._299_  (.A(\u_usb_host.u_core._062_ ),
    .B(\u_usb_host.u_core._114_ ),
    .Y(\u_usb_host.u_core._115_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core._300_  (.A1(\u_usb_host.u_core._062_ ),
    .A2(\u_usb_host.u_core._114_ ),
    .B1(\u_usb_host.u_core._115_ ),
    .C1(\u_usb_host.u_core._073_ ),
    .X(\u_usb_host.u_core._012_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_core._301_  (.A1(\u_usb_host.u_core.sof_time_q[13] ),
    .A2(\u_usb_host.u_core.sof_time_q[14] ),
    .A3(\u_usb_host.u_core._079_ ),
    .A4(\u_usb_host.u_core._109_ ),
    .B1(\u_usb_host.u_core.sof_time_q[15] ),
    .X(\u_usb_host.u_core._116_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core._302_  (.A1(\u_usb_host.u_core._067_ ),
    .A2(\u_usb_host.u_core._114_ ),
    .B1(\u_usb_host.u_core._116_ ),
    .C1(\u_usb_host.u_core._073_ ),
    .X(\u_usb_host.u_core._013_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._303_  (.A0(\u_usb_host.u_core._064_ ),
    .A1(\u_usb_host.u_core._086_ ),
    .S(\u_usb_host.u_core._002_ ),
    .X(\u_usb_host.u_core._023_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._304_  (.A(\u_usb_host.u_core.usb_xfer_token_in_out_w ),
    .B(\u_usb_host.u_core._073_ ),
    .X(\u_usb_host.u_core._049_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._305_  (.A(\u_usb_host.u_core.usb_xfer_token_ack_out_w ),
    .B(\u_usb_host.u_core._073_ ),
    .X(\u_usb_host.u_core._048_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._306_  (.A(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ),
    .X(\u_usb_host.u_core.token_pid_w[0] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._307_  (.A_N(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ),
    .X(\u_usb_host.u_core.token_pid_w[1] ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._308_  (.A(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ),
    .X(\u_usb_host.u_core.token_pid_w[2] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._309_  (.A_N(\u_usb_host.u_core.sof_transfer_q ),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ),
    .X(\u_usb_host.u_core.token_pid_w[3] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._310_  (.A_N(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ),
    .X(\u_usb_host.u_core.token_pid_w[4] ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._311_  (.A(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ),
    .X(\u_usb_host.u_core.token_pid_w[5] ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core._312_  (.A_N(\u_usb_host.u_core.sof_transfer_q ),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ),
    .X(\u_usb_host.u_core.token_pid_w[6] ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._313_  (.A(net525),
    .B(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ),
    .X(\u_usb_host.u_core.token_pid_w[7] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._314_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ),
    .A1(\u_usb_host.u_core.sof_value_q[6] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._315_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ),
    .A1(\u_usb_host.u_core.sof_value_q[5] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[1] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._316_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ),
    .A1(\u_usb_host.u_core.sof_value_q[4] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[2] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._317_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ),
    .A1(\u_usb_host.u_core.sof_value_q[3] ),
    .S(net525),
    .X(\u_usb_host.u_core.token_dev_w[3] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._318_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ),
    .A1(\u_usb_host.u_core.sof_value_q[2] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[4] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._319_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ),
    .A1(\u_usb_host.u_core.sof_value_q[1] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[5] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._320_  (.A0(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ),
    .A1(\u_usb_host.u_core.sof_value_q[0] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_dev_w[6] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._321_  (.A0(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ),
    .A1(\u_usb_host.u_core.sof_value_q[10] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_ep_w[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._322_  (.A0(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ),
    .A1(\u_usb_host.u_core.sof_value_q[9] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_ep_w[1] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._323_  (.A0(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ),
    .A1(\u_usb_host.u_core.sof_value_q[8] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_ep_w[2] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core._324_  (.A0(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ),
    .A1(\u_usb_host.u_core.sof_value_q[7] ),
    .S(net524),
    .X(\u_usb_host.u_core.token_ep_w[3] ));
 sky130_fd_sc_hd__nor3_2 \u_usb_host.u_core._325_  (.A(\u_usb_host.u_core._063_ ),
    .B(\u_usb_host.u_core._087_ ),
    .C(\u_usb_host.u_core._089_ ),
    .Y(\u_usb_host.u_core._117_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._326_  (.A1(\u_usb_host.u_core.usb_xfer_token_ack_out_w ),
    .A2(net96),
    .B1(net89),
    .B2(\u_usb_host.u_core.sof_time_q[13] ),
    .X(\u_usb_host.u_core._118_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._327_  (.A1(net578),
    .A2(net88),
    .B1(\u_usb_host.u_core._118_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[29] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._328_  (.A1(net588),
    .A2(net94),
    .B1(net89),
    .B2(\u_usb_host.u_core.sof_time_q[12] ),
    .X(\u_usb_host.u_core._119_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._329_  (.A1(net113),
    .A2(net87),
    .B1(\u_usb_host.u_core._119_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[28] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._330_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ),
    .A2(net96),
    .B1(net89),
    .B2(\u_usb_host.u_core.sof_time_q[0] ),
    .X(\u_usb_host.u_core._120_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._331_  (.A1(\u_usb_host.u_core.status_response_w[0] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._120_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[16] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._332_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ),
    .A2(net95),
    .B1(net89),
    .B2(\u_usb_host.u_core.sof_time_q[1] ),
    .X(\u_usb_host.u_core._121_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._333_  (.A1(\u_usb_host.u_core.status_response_w[1] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._121_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[17] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._334_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ),
    .A2(net95),
    .B1(net90),
    .B2(\u_usb_host.u_core.sof_time_q[2] ),
    .X(\u_usb_host.u_core._122_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._335_  (.A1(\u_usb_host.u_core.status_response_w[2] ),
    .A2(net87),
    .B1(\u_usb_host.u_core._122_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[18] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._336_  (.A1(\u_usb_host.u_core.sof_time_q[3] ),
    .A2(net90),
    .B1(net86),
    .B2(\u_usb_host.u_core.status_response_w[3] ),
    .X(\u_usb_host.u_core._123_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._337_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ),
    .A2(net95),
    .B1(\u_usb_host.u_core._123_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[19] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._338_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ),
    .A2(net94),
    .B1(net90),
    .B2(\u_usb_host.u_core.sof_time_q[4] ),
    .X(\u_usb_host.u_core._124_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._339_  (.A1(\u_usb_host.u_core.status_response_w[4] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._124_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[20] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._340_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ),
    .A2(net95),
    .B1(net90),
    .B2(\u_usb_host.u_core.sof_time_q[5] ),
    .X(\u_usb_host.u_core._125_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._341_  (.A1(\u_usb_host.u_core.status_response_w[5] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._125_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[21] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._342_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ),
    .A2(net94),
    .B1(net90),
    .B2(\u_usb_host.u_core.sof_time_q[6] ),
    .X(\u_usb_host.u_core._126_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._343_  (.A1(\u_usb_host.u_core.status_response_w[6] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._126_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[22] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._344_  (.A1(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ),
    .A2(net95),
    .B1(net90),
    .B2(\u_usb_host.u_core.sof_time_q[7] ),
    .X(\u_usb_host.u_core._127_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._345_  (.A1(\u_usb_host.u_core.status_response_w[7] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._127_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[23] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._346_  (.A1(\u_usb_host.u_core.utmi_xcvrselect_o[1] ),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(\u_usb_host.u_core._098_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.data_o[4] ),
    .X(\u_usb_host.u_core._128_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._347_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[4] ),
    .A2(net92),
    .B1(net88),
    .B2(\u_usb_host.u_core.status_rx_count_w[4] ),
    .X(\u_usb_host.u_core._129_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._348_  (.A(\u_usb_host.u_core._128_ ),
    .B(\u_usb_host.u_core._129_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[4] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._349_  (.A1(\u_usb_host.u_core.sof_time_q[15] ),
    .A2(net89),
    .B1(net87),
    .B2(net583),
    .X(\u_usb_host.u_core.reg_rdata_r[31] ));
 sky130_fd_sc_hd__nor3_2 \u_usb_host.u_core._350_  (.A(\u_usb_host.u_core._063_ ),
    .B(\u_usb_host.u_core._089_ ),
    .C(\u_usb_host.u_core._093_ ),
    .Y(\u_usb_host.u_core._130_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._351_  (.A1(net592),
    .A2(\u_usb_host.u_core._095_ ),
    .B1(\u_usb_host.u_core._130_ ),
    .B2(\u_usb_host.u_core.intr_sof_q ),
    .X(\u_usb_host.u_core._131_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._352_  (.A1(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[0] ),
    .X(\u_usb_host.u_core._132_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._353_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[0] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(net91),
    .B2(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .C1(\u_usb_host.u_core._132_ ),
    .X(\u_usb_host.u_core._133_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._354_  (.A1(\u_usb_host.u_core.status_rx_count_w[0] ),
    .A2(\u_usb_host.u_core._117_ ),
    .B1(net593),
    .C1(\u_usb_host.u_core._133_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[0] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._355_  (.A1(net612),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[6] ),
    .X(\u_usb_host.u_core._134_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._356_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ),
    .A2(net96),
    .B1(net88),
    .B2(\u_usb_host.u_core.status_rx_count_w[6] ),
    .X(\u_usb_host.u_core._135_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._357_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[6] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(\u_usb_host.u_core._134_ ),
    .C1(\u_usb_host.u_core._135_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[6] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._358_  (.A1(\u_usb_host.u_core.utmi_xcvrselect_o[0] ),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[3] ),
    .X(\u_usb_host.u_core._136_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._359_  (.A1(net589),
    .A2(\u_usb_host.u_core._095_ ),
    .B1(\u_usb_host.u_core._098_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.data_o[3] ),
    .X(\u_usb_host.u_core._137_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._360_  (.A1(\u_usb_host.u_core.status_rx_count_w[3] ),
    .A2(net88),
    .B1(\u_usb_host.u_core._136_ ),
    .C1(\u_usb_host.u_core._137_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[3] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._361_  (.A1(net594),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[5] ),
    .X(\u_usb_host.u_core._138_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._362_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ),
    .A2(net96),
    .B1(net88),
    .B2(\u_usb_host.u_core.status_rx_count_w[5] ),
    .X(\u_usb_host.u_core._139_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._363_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[5] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(\u_usb_host.u_core._138_ ),
    .C1(\u_usb_host.u_core._139_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[5] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._364_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[2] ),
    .A2(net93),
    .B1(net91),
    .B2(net585),
    .X(\u_usb_host.u_core._140_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._365_  (.A1(\u_usb_host.u_core.status_rx_count_w[2] ),
    .A2(net88),
    .B1(\u_usb_host.u_core._130_ ),
    .B2(\u_usb_host.u_core.intr_err_q ),
    .X(\u_usb_host.u_core._141_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._366_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[1] ),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(\u_usb_host.u_core._095_ ),
    .B2(\u_usb_host.u_core.usb_irq_mask_err_out_w ),
    .C1(\u_usb_host.u_core._141_ ),
    .X(\u_usb_host.u_core._142_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._367_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[2] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(\u_usb_host.u_core._140_ ),
    .C1(\u_usb_host.u_core._142_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[2] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._368_  (.A1(net601),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[7] ),
    .X(\u_usb_host.u_core._143_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._369_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ),
    .A2(net96),
    .B1(net88),
    .B2(\u_usb_host.u_core.status_rx_count_w[7] ),
    .X(\u_usb_host.u_core._144_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._370_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[7] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(\u_usb_host.u_core._143_ ),
    .C1(\u_usb_host.u_core._144_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[7] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._371_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[0] ),
    .A2(\u_usb_host.u_core._094_ ),
    .B1(\u_usb_host.u_core._130_ ),
    .B2(net590),
    .X(\u_usb_host.u_core._145_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._372_  (.A1(\u_usb_host.u_core.usb_irq_mask_done_out_w ),
    .A2(\u_usb_host.u_core._095_ ),
    .B1(net93),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[1] ),
    .X(\u_usb_host.u_core._146_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._373_  (.A1(\u_usb_host.u_core.u_fifo_rx.data_o[1] ),
    .A2(\u_usb_host.u_core._098_ ),
    .B1(net91),
    .B2(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .C1(\u_usb_host.u_core._146_ ),
    .X(\u_usb_host.u_core._147_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core._374_  (.A1(\u_usb_host.u_core.status_rx_count_w[1] ),
    .A2(net88),
    .B1(\u_usb_host.u_core._145_ ),
    .C1(\u_usb_host.u_core._147_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[1] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._375_  (.A1(\u_usb_host.u_core.usb_xfer_token_in_out_w ),
    .A2(net96),
    .B1(net89),
    .B2(\u_usb_host.u_core.sof_time_q[14] ),
    .X(\u_usb_host.u_core._148_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._376_  (.A1(net576),
    .A2(net87),
    .B1(\u_usb_host.u_core._148_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[30] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._377_  (.A1(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[8] ),
    .X(\u_usb_host.u_core._149_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._378_  (.A1(\u_usb_host.u_core.status_rx_count_w[8] ),
    .A2(net88),
    .B1(\u_usb_host.u_core._149_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[8] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._379_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[9] ),
    .X(\u_usb_host.u_core._150_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._380_  (.A1(\u_usb_host.u_core.status_rx_count_w[9] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._150_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[9] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._381_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[10] ),
    .X(\u_usb_host.u_core._151_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._382_  (.A1(\u_usb_host.u_core.status_rx_count_w[10] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._151_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[10] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._383_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ),
    .A2(net95),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[11] ),
    .X(\u_usb_host.u_core._152_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._384_  (.A1(\u_usb_host.u_core.status_rx_count_w[11] ),
    .A2(net86),
    .B1(\u_usb_host.u_core._152_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[11] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._385_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[12] ),
    .X(\u_usb_host.u_core._153_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._386_  (.A1(\u_usb_host.u_core.status_rx_count_w[12] ),
    .A2(net87),
    .B1(\u_usb_host.u_core._153_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[12] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._387_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[13] ),
    .X(\u_usb_host.u_core._154_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._388_  (.A1(\u_usb_host.u_core.status_rx_count_w[13] ),
    .A2(net87),
    .B1(\u_usb_host.u_core._154_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[13] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._389_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[14] ),
    .X(\u_usb_host.u_core._155_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._390_  (.A1(\u_usb_host.u_core.status_rx_count_w[14] ),
    .A2(net87),
    .B1(\u_usb_host.u_core._155_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[14] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._391_  (.A1(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ),
    .A2(net94),
    .B1(net92),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[15] ),
    .X(\u_usb_host.u_core._156_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core._392_  (.A1(\u_usb_host.u_core.status_rx_count_w[15] ),
    .A2(net87),
    .B1(\u_usb_host.u_core._156_ ),
    .X(\u_usb_host.u_core.reg_rdata_r[15] ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_core._393_  (.A(\u_usb_host.reg_ack ),
    .B(\u_usb_host.reg_wr ),
    .C_N(\u_usb_host.reg_cs ),
    .X(\u_usb_host.u_core._046_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_core._394_  (.A(\u_usb_host.u_core._046_ ),
    .Y(\u_usb_host.u_core._033_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._395_  (.A(\u_usb_host.reg_wdata[31] ),
    .B(\u_usb_host.u_core._037_ ),
    .X(\u_usb_host.u_core._032_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core._396_  (.A(\u_usb_host.u_core._090_ ),
    .B(\u_usb_host.u_core._093_ ),
    .Y(\u_usb_host.u_core._157_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._397_  (.A(\u_usb_host.reg_wdata[0] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._030_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._398_  (.A(\u_usb_host.reg_wdata[1] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._028_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._399_  (.A(\u_usb_host.reg_wdata[2] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._029_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._400_  (.A(\u_usb_host.reg_wdata[3] ),
    .B(\u_usb_host.u_core._157_ ),
    .X(\u_usb_host.u_core._027_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._401_  (.A(\u_usb_host.u_core.cfg_wr ),
    .B(\u_usb_host.reg_wdata[8] ),
    .C(\u_usb_host.u_core._094_ ),
    .X(\u_usb_host.u_core._024_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._402_  (.A(\u_usb_host.u_core._098_ ),
    .B(\u_usb_host.u_core._033_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.pop_i ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core._403_  (.A1(\u_usb_host.u_core.usb_irq_mask_done_out_w ),
    .A2(\u_usb_host.u_core.intr_done_q ),
    .B1(\u_usb_host.u_core.device_det_q ),
    .B2(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ),
    .X(\u_usb_host.u_core._158_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core._404_  (.A1(\u_usb_host.u_core.usb_irq_mask_sof_out_w ),
    .A2(\u_usb_host.u_core.intr_sof_q ),
    .B1(\u_usb_host.u_core.usb_irq_mask_err_out_w ),
    .B2(\u_usb_host.u_core.intr_err_q ),
    .C1(\u_usb_host.u_core._158_ ),
    .X(\u_usb_host.u_core._005_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._405_  (.A(\u_usb_host.u_core.sof_value_q[0] ),
    .B(\u_usb_host.u_core.sof_value_q[1] ),
    .X(\u_usb_host.u_core._052_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._406_  (.A(\u_usb_host.u_core.sof_value_q[0] ),
    .B(\u_usb_host.u_core.sof_value_q[2] ),
    .C(\u_usb_host.u_core.sof_value_q[1] ),
    .X(\u_usb_host.u_core._159_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._407_  (.A1(\u_usb_host.u_core.sof_value_q[0] ),
    .A2(\u_usb_host.u_core.sof_value_q[1] ),
    .B1(\u_usb_host.u_core.sof_value_q[2] ),
    .Y(\u_usb_host.u_core._160_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._408_  (.A(\u_usb_host.u_core._159_ ),
    .B(\u_usb_host.u_core._160_ ),
    .Y(\u_usb_host.u_core._053_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core._409_  (.A(\u_usb_host.u_core.sof_value_q[0] ),
    .B(\u_usb_host.u_core.sof_value_q[3] ),
    .C(\u_usb_host.u_core.sof_value_q[2] ),
    .D(\u_usb_host.u_core.sof_value_q[1] ),
    .X(\u_usb_host.u_core._161_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._410_  (.A(\u_usb_host.u_core.sof_value_q[3] ),
    .B(\u_usb_host.u_core._159_ ),
    .Y(\u_usb_host.u_core._162_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._411_  (.A(\u_usb_host.u_core._161_ ),
    .B(\u_usb_host.u_core._162_ ),
    .Y(\u_usb_host.u_core._054_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._412_  (.A(\u_usb_host.u_core.sof_value_q[4] ),
    .B(\u_usb_host.u_core._161_ ),
    .X(\u_usb_host.u_core._055_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._413_  (.A(\u_usb_host.u_core.sof_value_q[5] ),
    .B(\u_usb_host.u_core.sof_value_q[4] ),
    .C(\u_usb_host.u_core._161_ ),
    .X(\u_usb_host.u_core._163_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._414_  (.A1(\u_usb_host.u_core.sof_value_q[4] ),
    .A2(\u_usb_host.u_core._161_ ),
    .B1(\u_usb_host.u_core.sof_value_q[5] ),
    .Y(\u_usb_host.u_core._164_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._415_  (.A(\u_usb_host.u_core._163_ ),
    .B(\u_usb_host.u_core._164_ ),
    .Y(\u_usb_host.u_core._056_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._416_  (.A(\u_usb_host.u_core.sof_value_q[6] ),
    .B(\u_usb_host.u_core._163_ ),
    .X(\u_usb_host.u_core._165_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._417_  (.A(\u_usb_host.u_core.sof_value_q[6] ),
    .B(\u_usb_host.u_core._163_ ),
    .Y(\u_usb_host.u_core._166_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._418_  (.A(\u_usb_host.u_core._165_ ),
    .B(\u_usb_host.u_core._166_ ),
    .Y(\u_usb_host.u_core._057_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core._419_  (.A(\u_usb_host.u_core.sof_value_q[7] ),
    .B(\u_usb_host.u_core._165_ ),
    .X(\u_usb_host.u_core._058_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core._420_  (.A(\u_usb_host.u_core.sof_value_q[8] ),
    .B(\u_usb_host.u_core.sof_value_q[7] ),
    .C(\u_usb_host.u_core._165_ ),
    .X(\u_usb_host.u_core._167_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core._421_  (.A1(\u_usb_host.u_core.sof_value_q[7] ),
    .A2(\u_usb_host.u_core._165_ ),
    .B1(\u_usb_host.u_core.sof_value_q[8] ),
    .Y(\u_usb_host.u_core._168_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core._422_  (.A(\u_usb_host.u_core._167_ ),
    .B(\u_usb_host.u_core._168_ ),
    .Y(\u_usb_host.u_core._059_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core._423_  (.A(\u_usb_host.u_core.sof_value_q[9] ),
    .B(\u_usb_host.u_core._167_ ),
    .Y(\u_usb_host.u_core._169_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core._424_  (.A(\u_usb_host.u_core.sof_value_q[9] ),
    .B(\u_usb_host.u_core._167_ ),
    .X(\u_usb_host.u_core._170_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core._425_  (.A(\u_usb_host.u_core._169_ ),
    .B(\u_usb_host.u_core._170_ ),
    .X(\u_usb_host.u_core._060_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core._426_  (.A(\u_usb_host.u_core.sof_value_q[10] ),
    .B(\u_usb_host.u_core._169_ ),
    .Y(\u_usb_host.u_core._051_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._427_  (.CLK(\u_usb_host.u_core._189_ ),
    .D(\u_usb_host.u_core._049_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.in_transfer_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._428_  (.CLK(\u_usb_host.u_core._187_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.utmi_dppulldown_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._429_  (.CLK(\u_usb_host.u_core._190_ ),
    .D(\u_usb_host.u_core.send_sof_w ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.sof_transfer_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._430_  (.CLK(\u_usb_host.u_core._191_ ),
    .D(\u_usb_host.u_core._048_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.resp_expected_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._431_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._171_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.utmi_xcvrselect_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._432_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._171_ ),
    .D(\u_usb_host.reg_wdata[4] ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.utmi_xcvrselect_o[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._433_  (.CLK(\u_usb_host.u_core._177_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_irq_mask_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._434_  (.CLK(\u_usb_host.u_core._199_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.utmi_termselect_o ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._435_  (.CLK(\u_usb_host.u_core._201_ ),
    .D(\u_usb_host.u_core._047_ ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.cfg_wr ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._436_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._437_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._438_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._439_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._440_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[4] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._441_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._442_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._443_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._444_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[8] ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._445_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[9] ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._446_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[10] ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._447_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[11] ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._448_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[12] ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._449_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[13] ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._450_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[14] ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._451_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._178_ ),
    .D(\u_usb_host.reg_wdata[15] ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.u_sie.data_len_i[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._452_  (.CLK(\u_usb_host.u_core._202_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.utmi_dmpulldown_o ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._453_  (.CLK(\u_usb_host.u_core._188_ ),
    .D(\u_usb_host.u_core._002_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.fifo_flush_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._454_  (.CLK(\u_usb_host.u_core._179_ ),
    .D(\u_usb_host.u_core._032_ ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.usb_rx_stat_start_pend_in_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._455_  (.CLK(\u_usb_host.u_core._180_ ),
    .D(\u_usb_host.reg_wdata[30] ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.usb_xfer_token_in_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._456_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[0] ),
    .RESET_B(net381),
    .Q(\u_usb_host.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._457_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(net591),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._458_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(net586),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._459_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[3] ),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._460_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[4] ),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._461_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[5] ),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._462_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[6] ),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._463_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[7] ),
    .RESET_B(net388),
    .Q(\u_usb_host.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._464_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[8] ),
    .RESET_B(net381),
    .Q(\u_usb_host.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._465_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[9] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._466_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[10] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._467_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[11] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._468_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[12] ),
    .RESET_B(net379),
    .Q(\u_usb_host.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._469_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[13] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._470_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[14] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._471_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[15] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._472_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[16] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._473_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[17] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._474_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[18] ),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._475_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[19] ),
    .RESET_B(net379),
    .Q(\u_usb_host.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._476_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[20] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._477_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[21] ),
    .RESET_B(net379),
    .Q(\u_usb_host.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._478_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[22] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._479_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[23] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._480_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[24] ),
    .RESET_B(net379),
    .Q(\u_usb_host.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._481_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[25] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._482_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[26] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._483_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[27] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._484_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[28] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._485_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core._200_ ),
    .D(net579),
    .RESET_B(net381),
    .Q(\u_usb_host.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._486_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core._200_ ),
    .D(net577),
    .RESET_B(net380),
    .Q(\u_usb_host.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._487_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core._200_ ),
    .D(\u_usb_host.u_core.reg_rdata_r[31] ),
    .RESET_B(net378),
    .Q(\u_usb_host.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._488_  (.CLK(\u_usb_host.u_core._181_ ),
    .D(\u_usb_host.reg_wdata[29] ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.usb_xfer_token_ack_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._489_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._172_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net392),
    .Q(\u_usb_host.u_core.utmi_op_mode_o[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._490_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._172_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net388),
    .Q(\u_usb_host.u_core.utmi_op_mode_o[1] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._491_  (.CLK(\u_usb_host.u_core._182_ ),
    .D(\u_usb_host.reg_wdata[28] ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.u_sie.data_idx_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._492_  (.CLK(\u_usb_host.u_core._173_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_ctrl_enable_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._493_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[16] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._494_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[17] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._495_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[18] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._496_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[19] ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._497_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[20] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._498_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[21] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._499_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[22] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._500_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._183_ ),
    .D(\u_usb_host.reg_wdata[23] ),
    .RESET_B(net372),
    .Q(\u_usb_host.u_core.usb_xfer_token_pid_bits_out_w[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._501_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[9] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._502_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[10] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._503_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[11] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._504_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[12] ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._505_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[13] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._506_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[14] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._507_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._184_ ),
    .D(\u_usb_host.reg_wdata[15] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_dev_addr_out_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._508_  (.CLK(\u_usb_host.u_core._174_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_irq_mask_device_detect_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._509_  (.CLK(\u_usb_host.u_core._175_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_irq_mask_err_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._510_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._511_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._512_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._513_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._185_ ),
    .D(\u_usb_host.reg_wdata[8] ),
    .RESET_B(net371),
    .Q(\u_usb_host.u_core.usb_xfer_token_ep_addr_out_w[3] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._514_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[0] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._515_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._516_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[2] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._517_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[3] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[3] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._518_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[4] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._519_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[5] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._520_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[6] ),
    .RESET_B(net370),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._521_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._186_ ),
    .D(\u_usb_host.reg_wdata[7] ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.u_fifo_tx.data_i[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._522_  (.CLK(\u_usb_host.u_core._176_ ),
    .D(\u_usb_host.reg_wdata[1] ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_irq_mask_done_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._523_  (.CLK(\u_usb_host.u_core._198_ ),
    .D(\u_usb_host.u_core._000_ ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.device_det_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._524_  (.CLK(\u_usb_host.u_core._194_ ),
    .D(\u_usb_host.u_core._026_ ),
    .RESET_B(net416),
    .Q(\u_usb_host.u_core.usb_err_q ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._525_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._050_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._526_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._052_ ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.sof_value_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._527_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._053_ ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.sof_value_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._528_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._054_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.sof_value_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._529_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._055_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.sof_value_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._530_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._056_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.sof_value_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._531_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._057_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._532_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._058_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._533_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._059_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._534_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._060_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._535_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._192_ ),
    .D(\u_usb_host.u_core._051_ ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.sof_value_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._536_  (.CLK(\u_usb_host.u_core._195_ ),
    .D(\u_usb_host.u_core._003_ ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.intr_done_q ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core._537_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._007_ ),
    .RESET_B(net385),
    .Q(\u_usb_host.u_core.sof_time_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._538_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._014_ ),
    .RESET_B(net385),
    .Q(\u_usb_host.u_core.sof_time_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._539_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._015_ ),
    .RESET_B(net385),
    .Q(\u_usb_host.u_core.sof_time_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._540_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._016_ ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.sof_time_q[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._541_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._017_ ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.sof_time_q[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._542_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._018_ ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.sof_time_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._543_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._019_ ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.sof_time_q[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._544_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._020_ ),
    .RESET_B(net383),
    .Q(\u_usb_host.u_core.sof_time_q[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._545_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._021_ ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.sof_time_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._546_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._022_ ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.sof_time_q[9] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._547_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._008_ ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.sof_time_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._548_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._009_ ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.sof_time_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._549_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._010_ ),
    .RESET_B(net382),
    .Q(\u_usb_host.u_core.sof_time_q[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._550_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._011_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.sof_time_q[13] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core._551_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._012_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.sof_time_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._552_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core._193_ ),
    .D(\u_usb_host.u_core._013_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.sof_time_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._553_  (.CLK(\u_usb_host.u_core._196_ ),
    .D(net587),
    .RESET_B(net380),
    .Q(\u_usb_host.u_core.intr_sof_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._554_  (.CLK(\u_usb_host.u_core._197_ ),
    .D(\u_usb_host.u_core._004_ ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.intr_err_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._555_  (.CLK(clknet_leaf_1_usb_clk),
    .D(\u_usb_host.u_core._006_ ),
    .RESET_B(net366),
    .Q(\u_usb_host.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._556_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_core._025_ ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.usb_ctrl_wr_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._557_  (.CLK(clknet_leaf_4_usb_clk),
    .D(\u_usb_host.u_core._024_ ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.u_fifo_tx.flush_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._558_  (.CLK(clknet_leaf_9_usb_clk),
    .D(\u_usb_host.u_core._027_ ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_core.usb_irq_ack_device_detect_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._559_  (.CLK(clknet_leaf_8_usb_clk),
    .D(\u_usb_host.u_core._029_ ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.usb_irq_ack_err_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._560_  (.CLK(clknet_leaf_9_usb_clk),
    .D(\u_usb_host.u_core._028_ ),
    .RESET_B(net388),
    .Q(\u_usb_host.u_core.usb_irq_ack_done_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._561_  (.CLK(clknet_leaf_8_usb_clk),
    .D(\u_usb_host.u_core._030_ ),
    .RESET_B(net380),
    .Q(\u_usb_host.u_core.usb_irq_ack_sof_out_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._562_  (.CLK(clknet_leaf_4_usb_clk),
    .D(\u_usb_host.u_core._031_ ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.u_fifo_tx.push_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._563_  (.CLK(clknet_leaf_19_usb_clk),
    .D(\u_usb_host.u_core._023_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.transfer_start_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._564_  (.CLK(clknet_leaf_8_usb_clk),
    .D(\u_usb_host.u_core.send_sof_w ),
    .RESET_B(net381),
    .Q(\u_usb_host.u_core.sof_irq_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._565_  (.CLK(clknet_leaf_8_usb_clk),
    .D(\u_usb_host.u_core._001_ ),
    .RESET_B(net387),
    .Q(\u_usb_host.u_core.err_cond_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core._566_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_core._005_ ),
    .RESET_B(net389),
    .Q(net81));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._567_  (.CLK(clknet_leaf_12_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._171_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._568_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._172_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._569_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._173_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._570_  (.CLK(clknet_leaf_9_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._174_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._571_  (.CLK(clknet_leaf_9_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._175_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._572_  (.CLK(clknet_leaf_9_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._176_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._573_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._034_ ),
    .GCLK(\u_usb_host.u_core._177_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._574_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._035_ ),
    .GCLK(\u_usb_host.u_core._178_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._575_  (.CLK(clknet_leaf_5_usb_clk),
    .GATE(\u_usb_host.u_core._036_ ),
    .GCLK(\u_usb_host.u_core._179_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._576_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._180_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._577_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._181_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._578_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._182_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._579_  (.CLK(clknet_leaf_3_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._183_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._580_  (.CLK(clknet_leaf_6_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._184_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._581_  (.CLK(clknet_leaf_5_usb_clk),
    .GATE(\u_usb_host.u_core._037_ ),
    .GCLK(\u_usb_host.u_core._185_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_core._582_  (.CLK(clknet_leaf_5_usb_clk),
    .GATE(\u_usb_host.u_core.cfg_wr ),
    .GCLK(\u_usb_host.u_core._186_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._583_  (.CLK(clknet_leaf_14_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._187_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._584_  (.CLK(clknet_leaf_19_usb_clk),
    .GATE(\u_usb_host.u_core._038_ ),
    .GCLK(\u_usb_host.u_core._188_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._585_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core._039_ ),
    .GCLK(\u_usb_host.u_core._189_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._586_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core._039_ ),
    .GCLK(\u_usb_host.u_core._190_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._587_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core._039_ ),
    .GCLK(\u_usb_host.u_core._191_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._588_  (.CLK(clknet_leaf_6_usb_clk),
    .GATE(\u_usb_host.u_core.send_sof_w ),
    .GCLK(\u_usb_host.u_core._192_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core._589_  (.CLK(clknet_leaf_6_usb_clk),
    .GATE(\u_usb_host.u_core._040_ ),
    .GCLK(\u_usb_host.u_core._193_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._590_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_core._041_ ),
    .GCLK(\u_usb_host.u_core._194_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._591_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_core._042_ ),
    .GCLK(\u_usb_host.u_core._195_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._592_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._043_ ),
    .GCLK(\u_usb_host.u_core._196_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._593_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._044_ ),
    .GCLK(\u_usb_host.u_core._197_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._594_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_core._045_ ),
    .GCLK(\u_usb_host.u_core._198_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._595_  (.CLK(clknet_leaf_13_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._199_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_core._596_  (.CLK(clknet_leaf_8_usb_clk),
    .GATE(\u_usb_host.u_core._033_ ),
    .GCLK(\u_usb_host.u_core._200_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._597_  (.CLK(clknet_leaf_1_usb_clk),
    .GATE(\u_usb_host.u_core._046_ ),
    .GCLK(\u_usb_host.u_core._201_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core._598_  (.CLK(clknet_leaf_14_usb_clk),
    .GATE(\u_usb_host.u_core._025_ ),
    .GCLK(\u_usb_host.u_core._202_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_rx._0788_  (.A(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0443_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._0789_  (.A(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0444_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._0790_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0445_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_rx._0791_  (.A(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0446_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core.u_fifo_rx._0793_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0447_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_core.u_fifo_rx._0794_  (.A1(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B1(\u_usb_host.u_core.fifo_rx_push_w ),
    .X(\u_usb_host.u_core.u_fifo_rx._0448_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_fifo_rx._0795_  (.A1(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B1(\u_usb_host.u_core.fifo_rx_push_w ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0449_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0796_  (.A(net401),
    .B(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0450_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_rx._0797_  (.A(net401),
    .B(net443),
    .C(net442),
    .D(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0451_ ));
 sky130_fd_sc_hd__nand3b_4 \u_usb_host.u_core.u_fifo_rx._0798_  (.A_N(net444),
    .B(net447),
    .C(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0452_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0799_  (.A(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0039_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0800_  (.A(net444),
    .B(net446),
    .X(\u_usb_host.u_core.u_fifo_rx._0453_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_rx._0801_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .B(net441),
    .C(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0454_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_rx._0802_  (.A_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0455_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core.u_fifo_rx._0803_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0456_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0804_  (.A(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .B(net99),
    .Y(\u_usb_host.u_core.u_fifo_rx._0042_ ));
 sky130_fd_sc_hd__nand4b_4 \u_usb_host.u_core.u_fifo_rx._0805_  (.A_N(net443),
    .B(net441),
    .C(net445),
    .D(net446),
    .Y(\u_usb_host.u_core.u_fifo_rx._0457_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core.u_fifo_rx._0806_  (.A(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0458_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0807_  (.A(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .B(net98),
    .Y(\u_usb_host.u_core.u_fifo_rx._0037_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0808_  (.A(net444),
    .B(net446),
    .Y(\u_usb_host.u_core.u_fifo_rx._0459_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core.u_fifo_rx._0809_  (.A(net444),
    .B(net446),
    .C(net443),
    .X(\u_usb_host.u_core.u_fifo_rx._0460_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0810_  (.A(net442),
    .B(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0461_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0811_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0041_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_rx._0812_  (.A(net447),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .C(net441),
    .D_N(net445),
    .X(\u_usb_host.u_core.u_fifo_rx._0462_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0813_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0044_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_rx._0814_  (.A(net445),
    .B(net443),
    .C(net441),
    .D_N(net446),
    .X(\u_usb_host.u_core.u_fifo_rx._0463_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0815_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0043_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_rx._0816_  (.A(net443),
    .B(net441),
    .C_N(net444),
    .D_N(net446),
    .X(\u_usb_host.u_core.u_fifo_rx._0464_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0817_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0045_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0818_  (.A(net444),
    .B(net447),
    .C_N(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0465_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0819_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0054_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_rx._0820_  (.A(net447),
    .B(net441),
    .C_N(net443),
    .D_N(net444),
    .X(\u_usb_host.u_core.u_fifo_rx._0466_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0821_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0048_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0822_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0053_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_rx._0823_  (.A(net445),
    .B(net441),
    .C_N(net443),
    .D_N(net446),
    .X(\u_usb_host.u_core.u_fifo_rx._0467_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0824_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0047_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_rx._0825_  (.A(net447),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .C_N(net441),
    .D_N(net445),
    .X(\u_usb_host.u_core.u_fifo_rx._0468_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0826_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0052_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_rx._0827_  (.A(net444),
    .B(net443),
    .C_N(net441),
    .D_N(net446),
    .X(\u_usb_host.u_core.u_fifo_rx._0469_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0828_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0051_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_rx._0829_  (.A(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ),
    .C_N(net441),
    .X(\u_usb_host.u_core.u_fifo_rx._0470_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0830_  (.A(\u_usb_host.u_core.u_fifo_rx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0050_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_rx._0831_  (.A(net442),
    .B(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .D_N(net443),
    .X(\u_usb_host.u_core.u_fifo_rx._0471_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0832_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0046_ ));
 sky130_fd_sc_hd__nand2b_4 \u_usb_host.u_core.u_fifo_rx._0833_  (.A_N(net442),
    .B(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0472_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0834_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0049_ ));
 sky130_fd_sc_hd__nand3b_2 \u_usb_host.u_core.u_fifo_rx._0835_  (.A_N(net447),
    .B(\u_usb_host.u_core.u_fifo_rx._0451_ ),
    .C(net444),
    .Y(\u_usb_host.u_core.u_fifo_rx._0473_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0836_  (.A(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0040_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0837_  (.A(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0038_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0838_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0036_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0839_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0035_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0840_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0034_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0841_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0033_ ));
 sky130_fd_sc_hd__nand2b_4 \u_usb_host.u_core.u_fifo_rx._0842_  (.A_N(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0474_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0843_  (.A(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0062_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core.u_fifo_rx._0844_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0061_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core.u_fifo_rx._0845_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0475_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0846_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0060_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0847_  (.A(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0059_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0848_  (.A(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0058_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0849_  (.A(net99),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0057_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0850_  (.A(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0056_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0851_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0455_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0055_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0852_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0032_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0853_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0031_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0854_  (.A(\u_usb_host.u_core.u_fifo_rx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0030_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0855_  (.A(net98),
    .B(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0029_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0856_  (.A(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0028_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0857_  (.A(\u_usb_host.u_core.u_fifo_rx._0458_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0027_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0858_  (.A(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .B(net98),
    .Y(\u_usb_host.u_core.u_fifo_rx._0026_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_core.u_fifo_rx._0860_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.pop_i ),
    .X(\u_usb_host.u_core.u_fifo_rx._0476_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0861_  (.A(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0477_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0862_  (.A(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0478_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._0863_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0025_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0864_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0024_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0865_  (.A(\u_usb_host.u_core.fifo_flush_q ),
    .B(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0023_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0866_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0479_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0867_  (.A(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0022_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0868_  (.A(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0021_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0869_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0020_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0870_  (.A(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0480_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0871_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0480_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0019_ ));
 sky130_fd_sc_hd__or2_4 \u_usb_host.u_core.u_fifo_rx._0872_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0481_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0873_  (.A(\u_usb_host.u_core.u_fifo_rx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0076_ ));
 sky130_fd_sc_hd__nor3_2 \u_usb_host.u_core.u_fifo_rx._0874_  (.A(\u_usb_host.u_core.u_fifo_rx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0463_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0075_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0875_  (.A(\u_usb_host.u_core.u_fifo_rx._0454_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0074_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0876_  (.A(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0073_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0877_  (.A(\u_usb_host.u_core.u_fifo_rx._0473_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0072_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0878_  (.A(\u_usb_host.u_core.u_fifo_rx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0071_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0879_  (.A(\u_usb_host.u_core.u_fifo_rx._0465_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0070_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0880_  (.A(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0069_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0881_  (.A(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0068_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0882_  (.A(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0067_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0883_  (.A(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0066_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0884_  (.A(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0064_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0885_  (.A(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .B(net97),
    .Y(\u_usb_host.u_core.u_fifo_rx._0065_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0886_  (.A(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0475_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0063_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0887_  (.A(\u_usb_host.u_core.u_fifo_rx._0472_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0081_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0888_  (.A(\u_usb_host.u_core.u_fifo_rx._0471_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0078_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0889_  (.A(\u_usb_host.u_core.u_fifo_rx._0466_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0080_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0890_  (.A(\u_usb_host.u_core.u_fifo_rx._0467_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0079_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0891_  (.A(\u_usb_host.u_core.u_fifo_rx._0464_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0077_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0892_  (.A(\u_usb_host.u_core.u_fifo_rx._0468_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0084_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0893_  (.A(\u_usb_host.u_core.u_fifo_rx._0457_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0085_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0894_  (.A(\u_usb_host.u_core.u_fifo_rx._0470_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0082_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0895_  (.A(\u_usb_host.u_core.u_fifo_rx._0469_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0083_ ));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_core.u_fifo_rx._0896_  (.A1(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B1_N(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0000_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0897_  (.A(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0482_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_fifo_rx._0898_  (.A0(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .A1(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .S(\u_usb_host.u_core.u_fifo_rx._0482_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0001_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0899_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0483_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0900_  (.A(\u_usb_host.u_core.u_fifo_rx._0444_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0483_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0484_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_rx._0901_  (.A(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0485_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0902_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0486_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0903_  (.A1(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0485_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0486_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0484_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0002_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0904_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0444_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0487_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0905_  (.A(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0487_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0488_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_rx._0906_  (.A(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0489_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_rx._0907_  (.A(\u_usb_host.u_core.u_fifo_rx._0489_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0490_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._0908_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx.count[0] ),
    .A3(\u_usb_host.u_core.u_fifo_rx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0491_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0909_  (.A1(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0490_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0491_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0488_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0003_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0910_  (.A(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0492_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0911_  (.A(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0489_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0493_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0912_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0489_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0494_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_rx._0913_  (.A1_N(\u_usb_host.u_core.u_fifo_rx._0493_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_rx._0494_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0492_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0004_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0914_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0445_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0495_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0915_  (.A(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0495_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0496_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0916_  (.A(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_rx._0489_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0497_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0917_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0493_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0498_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_rx._0918_  (.A1_N(\u_usb_host.u_core.u_fifo_rx._0497_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_rx._0498_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0496_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0005_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_rx._0919_  (.A(\u_usb_host.u_core.u_fifo_rx._0443_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0497_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0499_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._0920_  (.A1(\u_usb_host.u_core.u_fifo_rx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0446_ ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0478_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0499_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0477_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0006_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_rx._0921_  (.A_N(net456),
    .B(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0007_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0922_  (.A(net456),
    .B(net453),
    .Y(\u_usb_host.u_core.u_fifo_rx._0500_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0923_  (.A(net456),
    .B(net453),
    .X(\u_usb_host.u_core.u_fifo_rx._0501_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0924_  (.A(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0500_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0501_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0008_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0925_  (.A1(net456),
    .A2(net453),
    .B1(net450),
    .X(\u_usb_host.u_core.u_fifo_rx._0502_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_rx._0926_  (.A(net456),
    .B(net453),
    .C(net450),
    .Y(\u_usb_host.u_core.u_fifo_rx._0503_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0927_  (.A(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0502_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0503_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0009_ ));
 sky130_fd_sc_hd__and4b_2 \u_usb_host.u_core.u_fifo_rx._0928_  (.A_N(net448),
    .B(net450),
    .C(net452),
    .D(net454),
    .X(\u_usb_host.u_core.u_fifo_rx._0504_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0929_  (.A(net448),
    .B(\u_usb_host.u_core.u_fifo_rx._0503_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0505_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_fifo_rx._0930_  (.A1(net363),
    .A2(\u_usb_host.u_core.u_fifo_rx._0505_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0010_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core.u_fifo_rx._0931_  (.A(net455),
    .B(net452),
    .C(net450),
    .D(net449),
    .X(\u_usb_host.u_core.u_fifo_rx._0506_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_rx._0932_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net362),
    .B1(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0507_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_fifo_rx._0933_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net362),
    .B1(\u_usb_host.u_core.u_fifo_rx._0507_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0011_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_rx._0934_  (.A_N(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0508_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_rx._0935_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0509_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_rx._0936_  (.A(net362),
    .B(net348),
    .Y(\u_usb_host.u_core.u_fifo_rx._0510_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0937_  (.A1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .A2(net362),
    .B1(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0511_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0938_  (.A(\u_usb_host.u_core.u_fifo_rx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0510_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0511_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0012_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0939_  (.A(net446),
    .B(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0013_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0940_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0453_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0459_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0014_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_rx._0941_  (.A1(net444),
    .A2(net446),
    .B1(net443),
    .X(\u_usb_host.u_core.u_fifo_rx._0512_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_core.u_fifo_rx._0942_  (.A_N(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0512_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0015_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_rx._0943_  (.A(net442),
    .B(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0513_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0944_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0513_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0016_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_fifo_rx._0945_  (.A(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0461_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0514_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_rx._0946_  (.A(\u_usb_host.u_core.u_fifo_rx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0514_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0017_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._0947_  (.A1(net442),
    .A2(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ),
    .A3(\u_usb_host.u_core.u_fifo_rx._0460_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0515_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0948_  (.A(\u_usb_host.u_core.u_fifo_rx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0480_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0515_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0018_ ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_core.u_fifo_rx._0949_  (.A(net454),
    .B(net453),
    .C(net451),
    .D(net449),
    .Y(\u_usb_host.u_core.u_fifo_rx._0516_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_rx._0950_  (.A(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0517_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0951_  (.A(net334),
    .B(net329),
    .X(\u_usb_host.u_core.u_fifo_rx._0518_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_rx._0952_  (.A(net334),
    .B(\u_usb_host.u_core.u_fifo_rx._0517_ ),
    .Y(\u_usb_host.u_core.u_fifo_rx._0519_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0953_  (.A_N(net453),
    .B_N(net450),
    .C(net448),
    .D(net454),
    .X(\u_usb_host.u_core.u_fifo_rx._0520_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0954_  (.A(net357),
    .B(net323),
    .X(\u_usb_host.u_core.u_fifo_rx._0521_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0955_  (.A(net455),
    .B(net450),
    .C(net448),
    .D_N(net452),
    .Y(\u_usb_host.u_core.u_fifo_rx._0522_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_rx._0956_  (.A_N(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0523_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0957_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][0] ),
    .B(net322),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0524_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0958_  (.A(net454),
    .B(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ),
    .C(net451),
    .D_N(net449),
    .Y(\u_usb_host.u_core.u_fifo_rx._0525_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0959_  (.A(net357),
    .B(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0526_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0960_  (.A_N(net454),
    .B_N(net450),
    .C(net448),
    .D(net453),
    .X(\u_usb_host.u_core.u_fifo_rx._0527_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0961_  (.A(net328),
    .B(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0528_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_rx._0962_  (.A_N(net451),
    .B(net449),
    .C(net455),
    .D(net452),
    .X(\u_usb_host.u_core.u_fifo_rx._0529_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0963_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][0] ),
    .B(net307),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0530_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_rx._0964_  (.A(net452),
    .B(net451),
    .C(net448),
    .D_N(net455),
    .Y(\u_usb_host.u_core.u_fifo_rx._0531_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0965_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][0] ),
    .B(net350),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0532_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0966_  (.A(net357),
    .B(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0533_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0967_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][0] ),
    .B(net343),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0534_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0968_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][0] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0535_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0969_  (.A(net329),
    .B(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0536_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0970_  (.A(net348),
    .B(\u_usb_host.u_core.u_fifo_rx._0525_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0537_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0971_  (.A(net329),
    .B(net323),
    .X(\u_usb_host.u_core.u_fifo_rx._0538_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0972_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][0] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0539_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0973_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][0] ),
    .B(net342),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0540_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0974_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][0] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0541_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0975_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][0] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0542_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0976_  (.A(net330),
    .B(\u_usb_host.u_core.u_fifo_rx._0522_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0543_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0977_  (.A_N(net450),
    .B_N(net448),
    .C(net455),
    .D(net452),
    .X(\u_usb_host.u_core.u_fifo_rx._0544_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0978_  (.A(net330),
    .B(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0545_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0979_  (.A(net358),
    .B(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0546_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0980_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][0] ),
    .B(net334),
    .C(net310),
    .X(\u_usb_host.u_core.u_fifo_rx._0547_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0981_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][0] ),
    .B(net313),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0548_ ));
 sky130_fd_sc_hd__nor4b_1 \u_usb_host.u_core.u_fifo_rx._0982_  (.A(net454),
    .B(net452),
    .C(net449),
    .D_N(net451),
    .Y(\u_usb_host.u_core.u_fifo_rx._0549_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0983_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][0] ),
    .B(net340),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0550_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0984_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][0] ),
    .B(net335),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0551_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0985_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][0] ),
    .B(net343),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0552_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0986_  (.A(net330),
    .B(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0553_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0987_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][0] ),
    .B(net340),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0554_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0988_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][0] ),
    .B(net330),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0555_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0989_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][0] ),
    .B(net337),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0556_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0990_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][0] ),
    .B(net314),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0557_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0991_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][0] ),
    .B(net316),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0558_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0992_  (.A(net357),
    .B(\u_usb_host.u_core.u_fifo_rx._0527_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0559_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0993_  (.A(net309),
    .B(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0560_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._0994_  (.A(net363),
    .B(net351),
    .X(\u_usb_host.u_core.u_fifo_rx._0561_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0995_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][0] ),
    .B(net362),
    .C(net342),
    .X(\u_usb_host.u_core.u_fifo_rx._0562_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._0996_  (.A_N(net454),
    .B_N(net453),
    .C(net451),
    .D(net449),
    .X(\u_usb_host.u_core.u_fifo_rx._0563_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0997_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][0] ),
    .B(net307),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0564_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._0998_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][0] ),
    .B(net314),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0565_ ));
 sky130_fd_sc_hd__and4b_2 \u_usb_host.u_core.u_fifo_rx._0999_  (.A_N(net452),
    .B(net451),
    .C(net449),
    .D(net455),
    .X(\u_usb_host.u_core.u_fifo_rx._0566_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1000_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][0] ),
    .B(net305),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0567_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1001_  (.A(net363),
    .B(net348),
    .X(\u_usb_host.u_core.u_fifo_rx._0568_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1002_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][0] ),
    .B(net359),
    .C(net305),
    .X(\u_usb_host.u_core.u_fifo_rx._0569_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1003_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][0] ),
    .B(net361),
    .C(net354),
    .X(\u_usb_host.u_core.u_fifo_rx._0570_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_rx._1004_  (.A_N(net453),
    .B_N(net448),
    .C(net450),
    .D(net454),
    .X(\u_usb_host.u_core.u_fifo_rx._0571_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1005_  (.A(net330),
    .B(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0572_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_rx._1006_  (.A_N(net454),
    .B(net452),
    .C(net451),
    .D(net448),
    .X(\u_usb_host.u_core.u_fifo_rx._0573_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1007_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][0] ),
    .B(net359),
    .C(net328),
    .X(\u_usb_host.u_core.u_fifo_rx._0574_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_rx._1008_  (.A_N(net454),
    .B_N(net448),
    .C(net450),
    .D(net452),
    .X(\u_usb_host.u_core.u_fifo_rx._0575_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1009_  (.A(net330),
    .B(\u_usb_host.u_core.u_fifo_rx._0575_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0576_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1010_  (.A(net330),
    .B(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0577_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1011_  (.A(net363),
    .B(net330),
    .X(\u_usb_host.u_core.u_fifo_rx._0578_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1012_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][0] ),
    .B(net343),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0579_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1013_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][0] ),
    .B(net306),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0580_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1014_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][0] ),
    .B(net363),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0581_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1015_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][0] ),
    .B(net354),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0582_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1016_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][0] ),
    .B(net343),
    .C(net285),
    .X(\u_usb_host.u_core.u_fifo_rx._0583_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1017_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][0] ),
    .B(net311),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0584_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1018_  (.A(net348),
    .B(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0585_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1019_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][0] ),
    .B(net354),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0586_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1020_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][0] ),
    .B(net340),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0587_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1021_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][0] ),
    .B(net325),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0588_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1022_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][0] ),
    .B(net355),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0589_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1023_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][0] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0590_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_rx._1024_  (.A(net358),
    .B(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0591_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1025_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][0] ),
    .B(net316),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0592_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1026_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0593_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1027_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[14][0] ),
    .A2(net327),
    .A3(net276),
    .B1(\u_usb_host.u_core.u_fifo_rx._0588_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0535_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0594_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1028_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0595_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1029_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0596_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1030_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0595_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0597_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1031_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0596_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0598_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1032_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][0] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0593_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0599_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1033_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][0] ),
    .A2(net355),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0589_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0600_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1034_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][0] ),
    .A2(net355),
    .A3(net279),
    .B1(\u_usb_host.u_core.u_fifo_rx._0600_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0547_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0601_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1035_  (.A(\u_usb_host.u_core.u_fifo_rx._0597_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0598_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0599_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0601_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0602_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1036_  (.A(\u_usb_host.u_core.u_fifo_rx._0551_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0567_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0569_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0580_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0603_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1037_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0564_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0530_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0541_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0604_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1038_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0542_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0539_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0532_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0605_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1039_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0586_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0582_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0570_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0606_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1040_  (.A(\u_usb_host.u_core.u_fifo_rx._0603_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0604_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0605_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0606_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0607_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1041_  (.A(\u_usb_host.u_core.u_fifo_rx._0540_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0555_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0562_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0590_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0608_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1042_  (.A(\u_usb_host.u_core.u_fifo_rx._0534_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0552_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0579_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0583_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0609_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1043_  (.A(\u_usb_host.u_core.u_fifo_rx._0524_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0548_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0557_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0565_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0610_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1044_  (.A(\u_usb_host.u_core.u_fifo_rx._0558_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0581_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0584_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0592_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0611_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1045_  (.A(\u_usb_host.u_core.u_fifo_rx._0608_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0609_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0610_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0611_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0612_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1046_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0613_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1047_  (.A(\u_usb_host.u_core.u_fifo_rx._0550_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0554_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0556_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0587_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0614_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1048_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0613_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0614_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0615_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1049_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0616_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1050_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][0] ),
    .A2(net328),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][0] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0617_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1051_  (.A(\u_usb_host.u_core.u_fifo_rx._0574_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0594_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0616_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0617_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0618_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1052_  (.A(\u_usb_host.u_core.u_fifo_rx._0607_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0612_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0615_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0618_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0619_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_rx._1053_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][0] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0602_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0619_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[0] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1054_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][1] ),
    .B(net316),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0620_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1055_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][1] ),
    .B(net315),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0621_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1056_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][1] ),
    .B(net308),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0622_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1057_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][1] ),
    .B(net349),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0623_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1058_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][1] ),
    .B(net343),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0624_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1059_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][1] ),
    .B(net315),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0625_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1060_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][1] ),
    .B(net337),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0626_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1061_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][1] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0627_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1062_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][1] ),
    .B(net347),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0628_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1063_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][1] ),
    .B(net335),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0629_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1064_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][1] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0630_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1065_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][1] ),
    .B(net334),
    .C(net319),
    .X(\u_usb_host.u_core.u_fifo_rx._0631_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1066_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][1] ),
    .B(net345),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0632_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1067_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][1] ),
    .B(net339),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0633_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1068_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][1] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0634_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1069_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][1] ),
    .B(net330),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0635_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1070_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][1] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0636_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1071_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][1] ),
    .B(net322),
    .C(net316),
    .X(\u_usb_host.u_core.u_fifo_rx._0637_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1072_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][1] ),
    .B(net362),
    .C(net338),
    .X(\u_usb_host.u_core.u_fifo_rx._0638_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1073_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][1] ),
    .B(net308),
    .C(net287),
    .X(\u_usb_host.u_core.u_fifo_rx._0639_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1074_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][1] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0640_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1075_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][1] ),
    .B(net354),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0641_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1076_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][1] ),
    .B(net311),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0642_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1077_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][1] ),
    .B(net325),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0643_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1078_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][1] ),
    .B(net359),
    .C(net329),
    .X(\u_usb_host.u_core.u_fifo_rx._0644_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1079_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][1] ),
    .B(net356),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0645_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1080_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][1] ),
    .B(net343),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0646_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1081_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][1] ),
    .B(net360),
    .C(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0647_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1082_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][1] ),
    .B(net360),
    .C(net351),
    .X(\u_usb_host.u_core.u_fifo_rx._0648_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1083_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][1] ),
    .B(net317),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0649_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1084_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][1] ),
    .B(net306),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0650_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1085_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][1] ),
    .B(net343),
    .C(net285),
    .X(\u_usb_host.u_core.u_fifo_rx._0651_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1086_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][1] ),
    .B(net304),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0652_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1087_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][1] ),
    .B(net339),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0653_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1088_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][1] ),
    .B(net339),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0654_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1089_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][1] ),
    .B(net351),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0655_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1090_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][1] ),
    .B(net315),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0656_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1091_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][1] ),
    .B(net363),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0657_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1092_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0658_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1093_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][1] ),
    .A2(net325),
    .A3(net283),
    .B1(\u_usb_host.u_core.u_fifo_rx._0634_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0643_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0659_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1094_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0660_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1095_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0661_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1096_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0660_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0662_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1097_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0661_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0663_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1098_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][1] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0658_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0664_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1099_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][1] ),
    .A2(net356),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0645_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0665_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1100_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][1] ),
    .A2(net356),
    .A3(net278),
    .B1(\u_usb_host.u_core.u_fifo_rx._0631_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0665_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0666_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1101_  (.A(\u_usb_host.u_core.u_fifo_rx._0662_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0663_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0664_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0666_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0667_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1102_  (.A(\u_usb_host.u_core.u_fifo_rx._0629_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0647_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0650_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0652_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0668_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1103_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0622_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0636_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0639_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0669_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1104_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0623_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0627_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0630_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0670_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1105_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0641_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0648_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0655_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0671_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1106_  (.A(\u_usb_host.u_core.u_fifo_rx._0668_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0669_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0670_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0671_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0672_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1107_  (.A(\u_usb_host.u_core.u_fifo_rx._0628_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0635_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0638_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0640_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0673_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1108_  (.A(\u_usb_host.u_core.u_fifo_rx._0624_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0632_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0646_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0651_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0674_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1109_  (.A(\u_usb_host.u_core.u_fifo_rx._0621_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0625_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0637_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0656_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0675_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1110_  (.A(\u_usb_host.u_core.u_fifo_rx._0620_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0642_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0649_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0657_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0676_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1111_  (.A(\u_usb_host.u_core.u_fifo_rx._0673_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0674_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0675_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0676_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0677_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1112_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0678_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1113_  (.A(\u_usb_host.u_core.u_fifo_rx._0626_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0633_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0653_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0654_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0679_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1114_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0678_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0679_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0680_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1115_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0681_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1116_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][1] ),
    .A2(net329),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][1] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0682_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1117_  (.A(\u_usb_host.u_core.u_fifo_rx._0644_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0659_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0681_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0682_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0683_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1118_  (.A(\u_usb_host.u_core.u_fifo_rx._0672_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0677_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0680_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0683_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0684_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1119_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][1] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0667_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0684_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[1] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1120_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][2] ),
    .B(net322),
    .C(net318),
    .X(\u_usb_host.u_core.u_fifo_rx._0685_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1121_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][2] ),
    .B(net308),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0686_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1122_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][2] ),
    .B(net349),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0687_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1123_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][2] ),
    .B(net319),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0688_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1124_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][2] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0689_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1125_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][2] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0690_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1126_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][2] ),
    .B(net342),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0691_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1127_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][2] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0692_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1128_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][2] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0693_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1129_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][2] ),
    .B(net334),
    .C(net310),
    .X(\u_usb_host.u_core.u_fifo_rx._0694_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1130_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][2] ),
    .B(net344),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0695_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1131_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][2] ),
    .B(net340),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0696_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1132_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][2] ),
    .B(net336),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0697_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1133_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][2] ),
    .B(net345),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0698_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1134_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][2] ),
    .B(net341),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0699_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1135_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][2] ),
    .B(net330),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0700_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1136_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][2] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0701_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1137_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][2] ),
    .B(net313),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0702_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1138_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][2] ),
    .B(net315),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0703_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1139_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][2] ),
    .B(net362),
    .C(net342),
    .X(\u_usb_host.u_core.u_fifo_rx._0704_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1140_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][2] ),
    .B(net307),
    .C(net287),
    .X(\u_usb_host.u_core.u_fifo_rx._0705_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1141_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][2] ),
    .B(net313),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0706_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1142_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][2] ),
    .B(net305),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0707_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1143_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][2] ),
    .B(net359),
    .C(net305),
    .X(\u_usb_host.u_core.u_fifo_rx._0708_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1144_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][2] ),
    .B(net360),
    .C(net351),
    .X(\u_usb_host.u_core.u_fifo_rx._0709_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1145_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][2] ),
    .B(net359),
    .C(net328),
    .X(\u_usb_host.u_core.u_fifo_rx._0710_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1146_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][2] ),
    .B(net344),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0711_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1147_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][2] ),
    .B(net306),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0712_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1148_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][2] ),
    .B(net363),
    .C(net312),
    .X(\u_usb_host.u_core.u_fifo_rx._0713_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1149_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][2] ),
    .B(net353),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0714_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1150_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][2] ),
    .B(net343),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0715_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1151_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][2] ),
    .B(net312),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0716_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1152_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][2] ),
    .B(net351),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0717_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1153_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][2] ),
    .B(net340),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0718_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1154_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][2] ),
    .B(net325),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0719_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1155_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][2] ),
    .B(net355),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0720_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1156_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][2] ),
    .B(net315),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0086_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1157_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][2] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0087_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1158_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0088_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1159_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[14][2] ),
    .A2(net325),
    .A3(net276),
    .B1(\u_usb_host.u_core.u_fifo_rx._0689_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0719_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0089_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1160_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0090_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1161_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0091_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1162_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0090_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0092_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1163_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0091_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0093_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1164_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][2] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0088_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0094_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1165_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][2] ),
    .A2(net355),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0720_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0095_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1166_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][2] ),
    .A2(net355),
    .A3(net279),
    .B1(\u_usb_host.u_core.u_fifo_rx._0694_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0095_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0096_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1167_  (.A(\u_usb_host.u_core.u_fifo_rx._0092_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0093_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0094_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0096_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0097_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1168_  (.A(\u_usb_host.u_core.u_fifo_rx._0697_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0707_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0708_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0712_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0098_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1169_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0686_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0692_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0705_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0099_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1170_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0687_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0690_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0693_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0100_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1171_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0709_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0714_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0717_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0101_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1172_  (.A(\u_usb_host.u_core.u_fifo_rx._0098_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0099_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0100_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0101_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0102_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1173_  (.A(\u_usb_host.u_core.u_fifo_rx._0691_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0700_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0704_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0087_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0103_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1174_  (.A(\u_usb_host.u_core.u_fifo_rx._0695_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0698_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0711_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0715_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0104_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1175_  (.A(\u_usb_host.u_core.u_fifo_rx._0685_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0688_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0702_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0706_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0105_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1176_  (.A(\u_usb_host.u_core.u_fifo_rx._0703_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0713_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0716_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0086_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0106_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1177_  (.A(\u_usb_host.u_core.u_fifo_rx._0103_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0104_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0105_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0106_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0107_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1178_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0108_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1179_  (.A(\u_usb_host.u_core.u_fifo_rx._0696_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0699_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0701_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0718_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0109_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1180_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0108_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0109_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0110_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1181_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0111_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1182_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][2] ),
    .A2(net328),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][2] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0112_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1183_  (.A(\u_usb_host.u_core.u_fifo_rx._0710_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0089_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0111_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0112_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0113_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1184_  (.A(\u_usb_host.u_core.u_fifo_rx._0102_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0107_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0110_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0113_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0114_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1185_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][2] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0097_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0114_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[2] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1186_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][3] ),
    .B(net314),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0115_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1187_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][3] ),
    .B(net308),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0116_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1188_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][3] ),
    .B(net349),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0117_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1189_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][3] ),
    .B(net314),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0118_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1190_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][3] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0119_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1191_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][3] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0120_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1192_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][3] ),
    .B(net342),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0121_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1193_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][3] ),
    .B(net323),
    .C(net310),
    .X(\u_usb_host.u_core.u_fifo_rx._0122_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1194_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][3] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0123_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1195_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][3] ),
    .B(net334),
    .C(net319),
    .X(\u_usb_host.u_core.u_fifo_rx._0124_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1196_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][3] ),
    .B(net344),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0125_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1197_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][3] ),
    .B(net340),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0126_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1198_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][3] ),
    .B(net336),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0127_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1199_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][3] ),
    .B(net344),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0128_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1200_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][3] ),
    .B(net340),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0129_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1201_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][3] ),
    .B(net331),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0130_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1202_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][3] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0131_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1203_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][3] ),
    .B(net322),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0132_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1204_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][3] ),
    .B(net311),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0133_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1205_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][3] ),
    .B(net362),
    .C(net338),
    .X(\u_usb_host.u_core.u_fifo_rx._0134_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1206_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][3] ),
    .B(net307),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0135_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1207_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][3] ),
    .B(net317),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0136_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1208_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][3] ),
    .B(net305),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0137_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1209_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][3] ),
    .B(net359),
    .C(net305),
    .X(\u_usb_host.u_core.u_fifo_rx._0138_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1210_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][3] ),
    .B(net360),
    .C(net351),
    .X(\u_usb_host.u_core.u_fifo_rx._0139_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1211_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][3] ),
    .B(net359),
    .C(net328),
    .X(\u_usb_host.u_core.u_fifo_rx._0140_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1212_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][3] ),
    .B(net356),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0141_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1213_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][3] ),
    .B(net344),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0142_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1214_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][3] ),
    .B(net306),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0143_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1215_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][3] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0144_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1216_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][3] ),
    .B(net353),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0145_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1217_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][3] ),
    .B(net344),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0146_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1218_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][3] ),
    .B(net311),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0147_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1219_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][3] ),
    .B(net351),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0148_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1220_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][3] ),
    .B(net314),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0149_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1221_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][3] ),
    .B(net340),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0150_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1222_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][3] ),
    .B(net325),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0151_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1223_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][3] ),
    .B(net363),
    .C(net311),
    .X(\u_usb_host.u_core.u_fifo_rx._0152_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1224_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0153_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1225_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[14][3] ),
    .A2(net327),
    .A3(net276),
    .B1(\u_usb_host.u_core.u_fifo_rx._0119_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0151_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0154_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1226_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0155_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1227_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0156_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1228_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0155_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0157_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1229_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0156_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0158_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1230_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][3] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0153_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0159_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1231_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][3] ),
    .A2(net356),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0141_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0160_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1232_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][3] ),
    .A2(net356),
    .A3(net278),
    .B1(\u_usb_host.u_core.u_fifo_rx._0124_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0160_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0161_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1233_  (.A(\u_usb_host.u_core.u_fifo_rx._0157_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0158_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0159_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0161_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0162_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1234_  (.A(\u_usb_host.u_core.u_fifo_rx._0127_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0137_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0138_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0143_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0163_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1235_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0116_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0122_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0135_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0164_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1236_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0117_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0120_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0123_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0165_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1237_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0139_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0145_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0148_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0166_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1238_  (.A(\u_usb_host.u_core.u_fifo_rx._0163_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0164_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0165_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0166_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0167_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1239_  (.A(\u_usb_host.u_core.u_fifo_rx._0121_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0130_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0134_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0144_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0168_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1240_  (.A(\u_usb_host.u_core.u_fifo_rx._0125_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0128_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0142_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0146_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0169_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1241_  (.A(\u_usb_host.u_core.u_fifo_rx._0115_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0118_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0132_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0149_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0170_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1242_  (.A(\u_usb_host.u_core.u_fifo_rx._0133_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0136_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0147_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0152_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0171_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1243_  (.A(\u_usb_host.u_core.u_fifo_rx._0168_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0169_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0170_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0171_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0172_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1244_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0173_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1245_  (.A(\u_usb_host.u_core.u_fifo_rx._0126_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0129_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0131_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0150_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0174_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1246_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0173_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0174_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0175_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1247_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0176_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1248_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][3] ),
    .A2(net328),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][3] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0177_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1249_  (.A(\u_usb_host.u_core.u_fifo_rx._0140_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0154_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0176_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0177_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0178_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1250_  (.A(\u_usb_host.u_core.u_fifo_rx._0167_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0172_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0175_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0178_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0179_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_rx._1251_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][3] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0162_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0179_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[3] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1252_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][4] ),
    .B(net352),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0180_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1253_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][4] ),
    .B(net322),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0181_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1254_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][4] ),
    .B(net345),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0182_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1255_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][4] ),
    .B(net308),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0183_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1256_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][4] ),
    .B(net331),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0184_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1257_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][4] ),
    .B(net315),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0185_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1258_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][4] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0186_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1259_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][4] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0187_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1260_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][4] ),
    .B(net342),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0188_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1261_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][4] ),
    .B(net334),
    .C(net310),
    .X(\u_usb_host.u_core.u_fifo_rx._0189_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1262_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][4] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0190_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1263_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][4] ),
    .B(net313),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0191_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1264_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][4] ),
    .B(net346),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0192_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1265_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][4] ),
    .B(net360),
    .C(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0193_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1266_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][4] ),
    .B(net341),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0194_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1267_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][4] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0195_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1268_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][4] ),
    .B(net336),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0196_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1269_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][4] ),
    .B(net313),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0197_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1270_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][4] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0198_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1271_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][4] ),
    .B(net313),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0199_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1272_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][4] ),
    .B(net362),
    .C(net342),
    .X(\u_usb_host.u_core.u_fifo_rx._0200_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1273_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][4] ),
    .B(net339),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0201_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1274_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][4] ),
    .B(net325),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0202_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1275_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][4] ),
    .B(net361),
    .C(net351),
    .X(\u_usb_host.u_core.u_fifo_rx._0203_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1276_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][4] ),
    .B(net326),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0204_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1277_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][4] ),
    .B(net307),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0205_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1278_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][4] ),
    .B(net359),
    .C(net326),
    .X(\u_usb_host.u_core.u_fifo_rx._0206_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1279_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0207_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1280_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][4] ),
    .B(net354),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0208_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1281_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][4] ),
    .B(net344),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0209_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1282_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][4] ),
    .B(net306),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0210_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1283_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][4] ),
    .B(net304),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0211_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1284_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][4] ),
    .B(net312),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0212_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1285_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][4] ),
    .B(net363),
    .C(net312),
    .X(\u_usb_host.u_core.u_fifo_rx._0213_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1286_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][4] ),
    .B(net346),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0214_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1287_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][4] ),
    .B(net339),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0215_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1288_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][4] ),
    .B(net338),
    .C(net279),
    .X(\u_usb_host.u_core.u_fifo_rx._0216_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1289_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][4] ),
    .B(net355),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0217_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1290_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][4] ),
    .B(net315),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0218_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1291_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][4] ),
    .B(net351),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0219_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1292_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0220_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1293_  (.A(\u_usb_host.u_core.u_fifo_rx._0195_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0202_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0204_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0206_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0221_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1294_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0222_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1295_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0207_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0223_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1296_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0222_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0224_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1297_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][4] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0220_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0225_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1298_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][4] ),
    .A2(net355),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0217_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0226_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1299_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][4] ),
    .A2(net355),
    .A3(net279),
    .B1(\u_usb_host.u_core.u_fifo_rx._0189_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0226_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0227_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1300_  (.A(\u_usb_host.u_core.u_fifo_rx._0223_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0224_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0225_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0227_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0228_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1301_  (.A(\u_usb_host.u_core.u_fifo_rx._0193_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0196_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0210_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0211_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0229_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1302_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0183_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0198_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0205_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0230_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1303_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0180_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0187_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0190_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0231_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1304_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0203_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0208_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0219_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0232_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1305_  (.A(\u_usb_host.u_core.u_fifo_rx._0229_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0230_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0231_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0232_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0233_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1306_  (.A(\u_usb_host.u_core.u_fifo_rx._0184_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0188_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0200_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0216_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0234_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1307_  (.A(\u_usb_host.u_core.u_fifo_rx._0182_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0192_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0209_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0214_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0235_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1308_  (.A(\u_usb_host.u_core.u_fifo_rx._0181_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0191_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0197_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0199_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0236_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1309_  (.A(\u_usb_host.u_core.u_fifo_rx._0185_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0212_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0213_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0218_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0237_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1310_  (.A(\u_usb_host.u_core.u_fifo_rx._0234_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0235_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0236_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0237_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0238_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1311_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0239_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1312_  (.A(\u_usb_host.u_core.u_fifo_rx._0186_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0194_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0201_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0215_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0240_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1313_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0239_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0240_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0241_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1314_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0242_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1315_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][4] ),
    .A2(net329),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][4] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0243_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._1316_  (.A(\u_usb_host.u_core.u_fifo_rx._0221_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0242_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0243_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0244_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1317_  (.A(\u_usb_host.u_core.u_fifo_rx._0233_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0238_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0241_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0244_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0245_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1318_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][4] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0228_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0245_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[4] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1319_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][5] ),
    .B(net322),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0246_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1320_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][5] ),
    .B(net345),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0247_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1321_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][5] ),
    .B(net307),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0248_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1322_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][5] ),
    .B(net331),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0249_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1323_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][5] ),
    .B(net311),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0250_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1324_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][5] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0251_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1325_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][5] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0252_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1326_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][5] ),
    .B(net347),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0253_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1327_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][5] ),
    .B(net336),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0254_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1328_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][5] ),
    .B(net352),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0255_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1329_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][5] ),
    .B(net352),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0256_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1330_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][5] ),
    .B(net313),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0257_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1331_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][5] ),
    .B(net345),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0258_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1332_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][5] ),
    .B(net304),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0259_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1333_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][5] ),
    .B(net339),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0260_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1334_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][5] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0261_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1335_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][5] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0262_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1336_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][5] ),
    .B(net313),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0263_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1337_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][5] ),
    .B(net334),
    .C(net319),
    .X(\u_usb_host.u_core.u_fifo_rx._0264_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1338_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][5] ),
    .B(net313),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0265_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1339_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][5] ),
    .B(net362),
    .C(net348),
    .X(\u_usb_host.u_core.u_fifo_rx._0266_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1340_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][5] ),
    .B(net353),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0267_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1341_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][5] ),
    .B(net325),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0268_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1342_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][5] ),
    .B(net309),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0269_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1343_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][5] ),
    .B(net327),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0270_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1344_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][5] ),
    .B(net359),
    .C(net326),
    .X(\u_usb_host.u_core.u_fifo_rx._0271_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1345_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0272_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1346_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][5] ),
    .B(net343),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0273_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1347_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][5] ),
    .B(net360),
    .C(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0274_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1348_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][5] ),
    .B(net360),
    .C(net353),
    .X(\u_usb_host.u_core.u_fifo_rx._0275_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1349_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][5] ),
    .B(net363),
    .C(net311),
    .X(\u_usb_host.u_core.u_fifo_rx._0276_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1350_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][5] ),
    .B(net345),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0277_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1351_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][5] ),
    .B(net305),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0278_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1352_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][5] ),
    .B(net312),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0279_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1353_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][5] ),
    .B(net339),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0280_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1354_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][5] ),
    .B(net338),
    .C(net279),
    .X(\u_usb_host.u_core.u_fifo_rx._0281_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1355_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][5] ),
    .B(net339),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0282_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1356_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][5] ),
    .B(net355),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0283_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1357_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][5] ),
    .B(net316),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0284_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1358_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][5] ),
    .B(net353),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0285_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1359_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0286_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1360_  (.A(\u_usb_host.u_core.u_fifo_rx._0261_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0268_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0270_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0271_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0287_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1361_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0288_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1362_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0272_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0289_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1363_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0288_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0290_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1364_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][5] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0286_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0291_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1365_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][5] ),
    .A2(net356),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0283_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0292_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1366_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][5] ),
    .A2(net356),
    .A3(net279),
    .B1(\u_usb_host.u_core.u_fifo_rx._0264_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0292_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0293_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1367_  (.A(\u_usb_host.u_core.u_fifo_rx._0289_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0290_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0291_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0293_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0294_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1368_  (.A(\u_usb_host.u_core.u_fifo_rx._0254_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0259_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0274_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0278_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0295_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1369_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0248_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0262_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0269_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0296_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1370_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0252_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0255_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0256_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0297_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1371_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0267_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0275_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0285_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0298_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1372_  (.A(\u_usb_host.u_core.u_fifo_rx._0295_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0296_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0297_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0298_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0299_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1373_  (.A(\u_usb_host.u_core.u_fifo_rx._0249_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0253_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0266_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0281_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0300_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1374_  (.A(\u_usb_host.u_core.u_fifo_rx._0247_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0258_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0273_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0277_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0301_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1375_  (.A(\u_usb_host.u_core.u_fifo_rx._0246_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0257_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0263_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0265_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0302_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1376_  (.A(\u_usb_host.u_core.u_fifo_rx._0250_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0276_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0279_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0284_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0303_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1377_  (.A(\u_usb_host.u_core.u_fifo_rx._0300_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0301_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0302_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0303_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0304_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1378_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0305_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1379_  (.A(\u_usb_host.u_core.u_fifo_rx._0251_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0260_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0280_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0282_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0306_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1380_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0305_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0306_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0307_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1381_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0308_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1382_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][5] ),
    .A2(net329),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][5] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0309_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._1383_  (.A(\u_usb_host.u_core.u_fifo_rx._0287_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0308_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0309_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0310_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1384_  (.A(\u_usb_host.u_core.u_fifo_rx._0299_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0304_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0307_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0310_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0311_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1385_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][5] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0294_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0311_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[5] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1386_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][6] ),
    .B(net322),
    .C(net318),
    .X(\u_usb_host.u_core.u_fifo_rx._0312_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1387_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][6] ),
    .B(net345),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0313_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1388_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][6] ),
    .B(net307),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0314_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1389_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][6] ),
    .B(net346),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0315_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1390_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][6] ),
    .B(net316),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0316_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1391_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][6] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0317_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1392_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][6] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0318_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1393_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][6] ),
    .B(net347),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0319_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1394_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][6] ),
    .B(net336),
    .C(net333),
    .X(\u_usb_host.u_core.u_fifo_rx._0320_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1395_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][6] ),
    .B(net352),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0321_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1396_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][6] ),
    .B(net351),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0322_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1397_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][6] ),
    .B(net314),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0323_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1398_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][6] ),
    .B(net331),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0324_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1399_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][6] ),
    .B(net306),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0325_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1400_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][6] ),
    .B(net341),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0326_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1401_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][6] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0327_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1402_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][6] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0328_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1403_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][6] ),
    .B(net313),
    .C(net298),
    .X(\u_usb_host.u_core.u_fifo_rx._0329_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1404_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][6] ),
    .B(net334),
    .C(net319),
    .X(\u_usb_host.u_core.u_fifo_rx._0330_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1405_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][6] ),
    .B(net314),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0331_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1406_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][6] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0506_ ),
    .C(net342),
    .X(\u_usb_host.u_core.u_fifo_rx._0332_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1407_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][6] ),
    .B(net353),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0333_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1408_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[13][6] ),
    .B(net326),
    .C(net283),
    .X(\u_usb_host.u_core.u_fifo_rx._0334_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1409_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][6] ),
    .B(net307),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0335_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1410_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][6] ),
    .B(net327),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0336_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1411_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][6] ),
    .B(net359),
    .C(net326),
    .X(\u_usb_host.u_core.u_fifo_rx._0337_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1412_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0338_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1413_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][6] ),
    .B(net344),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0339_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1414_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][6] ),
    .B(net360),
    .C(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0340_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1415_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][6] ),
    .B(net360),
    .C(net353),
    .X(\u_usb_host.u_core.u_fifo_rx._0341_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1416_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][6] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0504_ ),
    .C(net316),
    .X(\u_usb_host.u_core.u_fifo_rx._0342_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1417_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][6] ),
    .B(net346),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0343_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1418_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][6] ),
    .B(net304),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0344_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1419_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][6] ),
    .B(net311),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0345_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1420_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][6] ),
    .B(net341),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0346_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1421_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][6] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0347_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1422_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][6] ),
    .B(net339),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0348_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1423_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][6] ),
    .B(net357),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0349_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1424_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][6] ),
    .B(net316),
    .C(\u_usb_host.u_core.u_fifo_rx._0571_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0350_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1425_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][6] ),
    .B(net353),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0351_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1426_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0352_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1427_  (.A(\u_usb_host.u_core.u_fifo_rx._0327_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0334_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0336_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0337_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0353_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1428_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0354_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1429_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0338_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0355_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1430_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0354_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0356_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1431_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][6] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0352_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0357_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1432_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][6] ),
    .A2(net357),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0349_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0358_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1433_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][6] ),
    .A2(net357),
    .A3(net278),
    .B1(\u_usb_host.u_core.u_fifo_rx._0330_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0358_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0359_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1434_  (.A(\u_usb_host.u_core.u_fifo_rx._0355_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0356_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0357_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0359_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0360_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1435_  (.A(\u_usb_host.u_core.u_fifo_rx._0320_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0325_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0340_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0344_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0361_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1436_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0314_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0328_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0335_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0362_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1437_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0318_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0321_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0322_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0363_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1438_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0333_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0341_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0351_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0364_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1439_  (.A(\u_usb_host.u_core.u_fifo_rx._0361_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0362_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0363_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0364_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0365_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1440_  (.A(\u_usb_host.u_core.u_fifo_rx._0319_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0324_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0332_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0347_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0366_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1441_  (.A(\u_usb_host.u_core.u_fifo_rx._0313_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0315_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0339_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0343_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0367_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1442_  (.A(\u_usb_host.u_core.u_fifo_rx._0312_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0323_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0329_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0331_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0368_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1443_  (.A(\u_usb_host.u_core.u_fifo_rx._0316_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0342_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0345_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0350_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0369_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1444_  (.A(\u_usb_host.u_core.u_fifo_rx._0366_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0367_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0368_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0369_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0370_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1445_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0371_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1446_  (.A(\u_usb_host.u_core.u_fifo_rx._0317_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0326_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0346_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0348_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0372_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1447_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0371_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0372_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0373_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1448_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0374_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1449_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][6] ),
    .A2(net329),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][6] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0375_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_rx._1450_  (.A(\u_usb_host.u_core.u_fifo_rx._0353_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0374_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0375_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0376_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1451_  (.A(\u_usb_host.u_core.u_fifo_rx._0365_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0370_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0373_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0376_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0377_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1452_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][6] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0360_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0377_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[6] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1453_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[34][7] ),
    .B(net322),
    .C(net317),
    .X(\u_usb_host.u_core.u_fifo_rx._0378_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1454_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[58][7] ),
    .B(net345),
    .C(net301),
    .X(\u_usb_host.u_core.u_fifo_rx._0379_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1455_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[43][7] ),
    .B(net307),
    .C(net299),
    .X(\u_usb_host.u_core.u_fifo_rx._0380_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1456_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[8][7] ),
    .B(net331),
    .C(net302),
    .X(\u_usb_host.u_core.u_fifo_rx._0381_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1457_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[40][7] ),
    .B(net316),
    .C(net303),
    .X(\u_usb_host.u_core.u_fifo_rx._0382_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1458_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[50][7] ),
    .B(net337),
    .C(net321),
    .X(\u_usb_host.u_core.u_fifo_rx._0383_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1459_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[16][7] ),
    .B(net350),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0384_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1460_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[57][7] ),
    .B(net342),
    .C(net324),
    .X(\u_usb_host.u_core.u_fifo_rx._0385_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1461_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[48][7] ),
    .B(net336),
    .C(net332),
    .X(\u_usb_host.u_core.u_fifo_rx._0386_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1462_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[18][7] ),
    .B(net349),
    .C(net320),
    .X(\u_usb_host.u_core.u_fifo_rx._0387_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1463_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[17][7] ),
    .B(net349),
    .C(net297),
    .X(\u_usb_host.u_core.u_fifo_rx._0388_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1464_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[35][7] ),
    .B(net315),
    .C(net295),
    .X(\u_usb_host.u_core.u_fifo_rx._0389_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1465_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[59][7] ),
    .B(net345),
    .C(net300),
    .X(\u_usb_host.u_core.u_fifo_rx._0390_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1466_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[46][7] ),
    .B(net306),
    .C(net277),
    .X(\u_usb_host.u_core.u_fifo_rx._0391_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1467_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[51][7] ),
    .B(net340),
    .C(net294),
    .X(\u_usb_host.u_core.u_fifo_rx._0392_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1468_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[49][7] ),
    .B(net335),
    .C(net296),
    .X(\u_usb_host.u_core.u_fifo_rx._0393_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1469_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[41][7] ),
    .B(net323),
    .C(net309),
    .X(\u_usb_host.u_core.u_fifo_rx._0394_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1470_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[33][7] ),
    .B(net315),
    .C(\u_usb_host.u_core.u_fifo_rx._0531_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0395_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1471_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[32][7] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0516_ ),
    .C(net319),
    .X(\u_usb_host.u_core.u_fifo_rx._0396_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1472_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[63][7] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0506_ ),
    .C(net342),
    .X(\u_usb_host.u_core.u_fifo_rx._0397_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1473_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[36][7] ),
    .B(net315),
    .C(net293),
    .X(\u_usb_host.u_core.u_fifo_rx._0398_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1474_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[37][7] ),
    .B(net316),
    .C(net282),
    .X(\u_usb_host.u_core.u_fifo_rx._0399_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1475_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[20][7] ),
    .B(net353),
    .C(net291),
    .X(\u_usb_host.u_core.u_fifo_rx._0400_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1476_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[14][7] ),
    .B(net325),
    .C(net276),
    .X(\u_usb_host.u_core.u_fifo_rx._0401_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1477_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[15][7] ),
    .B(net361),
    .C(net328),
    .X(\u_usb_host.u_core.u_fifo_rx._0402_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1478_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[28][7] ),
    .B(net357),
    .C(net289),
    .X(\u_usb_host.u_core.u_fifo_rx._0403_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1479_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[60][7] ),
    .B(net343),
    .C(net290),
    .X(\u_usb_host.u_core.u_fifo_rx._0404_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1480_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[47][7] ),
    .B(net360),
    .C(net304),
    .X(\u_usb_host.u_core.u_fifo_rx._0405_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1481_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[31][7] ),
    .B(net361),
    .C(net354),
    .X(\u_usb_host.u_core.u_fifo_rx._0406_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1482_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[61][7] ),
    .B(net345),
    .C(net286),
    .X(\u_usb_host.u_core.u_fifo_rx._0407_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1483_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[45][7] ),
    .B(net304),
    .C(net284),
    .X(\u_usb_host.u_core.u_fifo_rx._0408_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1484_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[38][7] ),
    .B(net311),
    .C(net275),
    .X(\u_usb_host.u_core.u_fifo_rx._0409_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1485_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[62][7] ),
    .B(net338),
    .C(net278),
    .X(\u_usb_host.u_core.u_fifo_rx._0410_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1486_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[52][7] ),
    .B(net340),
    .C(net292),
    .X(\u_usb_host.u_core.u_fifo_rx._0411_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1487_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[39][7] ),
    .B(\u_usb_host.u_core.u_fifo_rx._0504_ ),
    .C(net311),
    .X(\u_usb_host.u_core.u_fifo_rx._0412_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1488_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[53][7] ),
    .B(net339),
    .C(net281),
    .X(\u_usb_host.u_core.u_fifo_rx._0413_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1489_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[44][7] ),
    .B(net307),
    .C(net288),
    .X(\u_usb_host.u_core.u_fifo_rx._0414_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_rx._1490_  (.A(\u_usb_host.u_core.u_fifo_rx.ram[21][7] ),
    .B(net353),
    .C(net280),
    .X(\u_usb_host.u_core.u_fifo_rx._0415_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1491_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[19][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[26][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0416_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1492_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[13][7] ),
    .A2(net325),
    .A3(net283),
    .B1(\u_usb_host.u_core.u_fifo_rx._0393_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0401_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0417_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1493_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[5][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[6][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0418_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1494_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[3][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[1][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0419_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1495_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[27][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[4][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0418_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0420_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1496_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[2][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[7][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0419_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0421_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_rx._1497_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[25][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[24][7] ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0416_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0422_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_rx._1498_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[29][7] ),
    .A2(net357),
    .A3(net285),
    .B1(\u_usb_host.u_core.u_fifo_rx._0403_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0423_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_rx._1499_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[30][7] ),
    .A2(net357),
    .A3(net278),
    .B1(\u_usb_host.u_core.u_fifo_rx._0396_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0423_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0424_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1500_  (.A(\u_usb_host.u_core.u_fifo_rx._0420_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0421_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0422_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0424_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0425_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1501_  (.A(\u_usb_host.u_core.u_fifo_rx._0386_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0391_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0405_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0408_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0426_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1502_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[42][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0380_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0394_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0414_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0427_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1503_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[23][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0384_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0387_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0388_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0428_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1504_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[22][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0400_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0406_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0415_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0429_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1505_  (.A(\u_usb_host.u_core.u_fifo_rx._0426_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0427_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0428_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0429_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0430_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1506_  (.A(\u_usb_host.u_core.u_fifo_rx._0381_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0385_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0397_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0410_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0431_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1507_  (.A(\u_usb_host.u_core.u_fifo_rx._0379_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0390_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0404_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0407_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0432_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1508_  (.A(\u_usb_host.u_core.u_fifo_rx._0378_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0389_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0395_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0398_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0433_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1509_  (.A(\u_usb_host.u_core.u_fifo_rx._0382_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0399_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0409_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0412_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0434_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1510_  (.A(\u_usb_host.u_core.u_fifo_rx._0431_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0432_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0433_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0434_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0435_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1511_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[55][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[54][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0436_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_rx._1512_  (.A(\u_usb_host.u_core.u_fifo_rx._0383_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0392_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0411_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0413_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0437_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_rx._1513_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[56][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0436_ ),
    .C1(\u_usb_host.u_core.u_fifo_rx._0437_ ),
    .D1(\u_usb_host.u_core.u_fifo_rx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0438_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_rx._1514_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[10][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[9][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0439_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_rx._1515_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[12][7] ),
    .A2(net328),
    .A3(net287),
    .B1(\u_usb_host.u_core.u_fifo_rx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx.ram[11][7] ),
    .X(\u_usb_host.u_core.u_fifo_rx._0440_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1516_  (.A(\u_usb_host.u_core.u_fifo_rx._0402_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0417_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0439_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0440_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0441_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_rx._1517_  (.A(\u_usb_host.u_core.u_fifo_rx._0430_ ),
    .B(\u_usb_host.u_core.u_fifo_rx._0435_ ),
    .C(\u_usb_host.u_core.u_fifo_rx._0438_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0441_ ),
    .X(\u_usb_host.u_core.u_fifo_rx._0442_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_fifo_rx._1518_  (.A1(\u_usb_host.u_core.u_fifo_rx.ram[0][7] ),
    .A2(\u_usb_host.u_core.u_fifo_rx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_rx._0425_ ),
    .B2(\u_usb_host.u_core.u_fifo_rx._0442_ ),
    .X(\u_usb_host.u_core.u_fifo_rx.data_o[7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1519_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1520_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1521_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1522_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1523_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1524_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1525_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1526_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0752_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1527_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1528_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net170),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1529_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1530_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1531_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1532_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1533_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1534_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0783_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1535_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1536_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1537_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1538_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1539_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1540_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1541_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1542_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0751_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1543_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1544_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1545_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1546_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1547_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1548_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1549_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1550_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0750_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1551_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1552_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net170),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1553_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1554_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1555_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1556_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(\u_usb_host.u_core.fifo_rx_data_w[5] ),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1557_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1558_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0782_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1559_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1560_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1561_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1562_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1563_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1564_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1565_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1566_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0749_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1567_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1568_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1569_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1570_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1571_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1572_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1573_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1574_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0781_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1575_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1576_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1577_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1578_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1579_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1580_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1581_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1582_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0748_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1583_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1584_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1585_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1586_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1587_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1588_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1589_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1590_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0747_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1591_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1592_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net170),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1593_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1594_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1595_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1596_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1597_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1598_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0780_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1599_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1600_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1601_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1602_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1603_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1604_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1605_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1606_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0746_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1607_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1608_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net170),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1609_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1610_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1611_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1612_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1613_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1614_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0779_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1615_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1616_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1617_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1618_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1619_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1620_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1621_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1622_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0745_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1623_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1624_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1625_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1626_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1627_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1628_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1629_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1630_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0744_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1631_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1632_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1633_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1634_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1635_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1636_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1637_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1638_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0778_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1639_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1640_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1641_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1642_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1643_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1644_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1645_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1646_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0743_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1647_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1648_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1649_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1650_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1651_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1652_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1653_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1654_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0777_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1655_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1656_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1657_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1658_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1659_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1660_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1661_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1662_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0742_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1663_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1664_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1665_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1666_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1667_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1668_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1669_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1670_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0741_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1671_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1672_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1673_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1674_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1675_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1676_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1677_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1678_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0776_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1679_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1680_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1681_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1682_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1683_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1684_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1685_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1686_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0740_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1687_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1688_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1689_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1690_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1691_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1692_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1693_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1694_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0775_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1695_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1696_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1697_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1698_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1699_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1700_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1701_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1702_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0739_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1703_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1704_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1705_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1706_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1707_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1708_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1709_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1710_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0738_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1711_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1712_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1713_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1714_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1715_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1716_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1717_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1718_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0774_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1719_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1720_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1721_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1722_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1723_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1724_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1725_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net134),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1726_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0737_ ),
    .D(net121),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1727_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net175),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1728_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1729_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net159),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1730_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net151),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1731_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net143),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1732_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net137),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1733_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net127),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1734_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0773_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1735_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1736_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1737_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1738_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1739_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1740_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1741_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1742_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0736_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1743_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1744_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1745_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1746_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1747_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1748_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1749_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1750_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0735_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1751_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1752_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1753_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1754_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1755_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1756_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1757_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1758_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0772_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1759_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1760_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1761_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1762_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1763_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1764_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1765_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1766_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0734_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1767_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1768_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1769_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net161),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1770_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1771_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1772_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net136),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1773_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1774_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0771_ ),
    .D(net119),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1775_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1776_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1777_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1778_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1779_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1780_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1781_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1782_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0733_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1783_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1784_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1785_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1786_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1787_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1788_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1789_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1790_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0732_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1791_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1792_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net168),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1793_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1794_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1795_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1796_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1797_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1798_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0770_ ),
    .D(net118),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1799_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1800_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1801_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1802_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1803_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1804_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1805_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1806_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0731_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1807_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1808_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1809_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1810_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1811_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1812_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1813_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1814_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0730_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1815_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1816_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net169),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1817_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1818_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net153),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1819_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1820_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1821_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1822_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0769_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1823_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1824_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1825_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1826_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1827_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1828_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1829_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1830_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0729_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1831_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1832_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1833_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1834_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1835_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1836_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1837_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1838_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0768_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1839_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1840_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1841_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1842_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1843_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1844_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1845_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1846_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0728_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1847_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1848_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net174),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1849_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1850_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1851_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1852_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1853_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1854_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0767_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[39][7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._1855_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0000_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._1856_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0001_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1857_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0002_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1858_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0003_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1859_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0004_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1860_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0005_ ),
    .RESET_B(net414),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1861_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0006_ ),
    .RESET_B(net411),
    .Q(\u_usb_host.u_core.u_fifo_rx.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1862_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1863_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1864_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1865_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1866_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1867_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1868_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1869_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0766_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[38][7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1870_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0007_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1871_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0008_ ),
    .RESET_B(net403),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1872_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0009_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1873_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0010_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._1874_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0011_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._1875_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0012_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_fifo_rx.rd_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1876_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1877_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1878_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1879_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1880_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1881_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1882_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1883_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0765_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1884_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1885_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1886_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1887_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1888_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1889_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1890_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1891_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0721_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1892_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1893_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1894_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1895_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1896_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1897_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1898_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1899_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0764_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1900_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1901_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1902_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1903_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1904_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1905_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1906_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1907_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0763_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[35][7] ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1908_  (.CLK(clknet_leaf_29_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0019_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0721_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1909_  (.CLK(clknet_leaf_29_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0020_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0722_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1910_  (.CLK(clknet_leaf_30_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0021_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0723_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1911_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0022_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0724_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1912_  (.CLK(clknet_leaf_21_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0023_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0725_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1913_  (.CLK(clknet_leaf_21_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0024_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0726_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1914_  (.CLK(clknet_leaf_23_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0025_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0727_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1915_  (.CLK(clknet_leaf_25_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0026_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0728_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1916_  (.CLK(clknet_leaf_23_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0027_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0729_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1917_  (.CLK(clknet_leaf_24_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0028_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0730_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1918_  (.CLK(clknet_leaf_23_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0029_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0731_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1919_  (.CLK(clknet_leaf_22_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0030_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0732_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1920_  (.CLK(clknet_leaf_22_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0031_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0733_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1921_  (.CLK(clknet_leaf_23_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0032_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0734_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1922_  (.CLK(clknet_leaf_24_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0033_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0735_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1923_  (.CLK(clknet_leaf_26_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0034_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0736_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1924_  (.CLK(clknet_leaf_20_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0035_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0737_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1925_  (.CLK(clknet_leaf_21_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0036_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0738_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1926_  (.CLK(clknet_leaf_36_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0037_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0739_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1927_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0038_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0740_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1928_  (.CLK(clknet_leaf_36_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0039_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0741_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1929_  (.CLK(clknet_leaf_36_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0040_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0742_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1930_  (.CLK(clknet_leaf_36_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0041_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0743_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1931_  (.CLK(clknet_leaf_40_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0042_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0744_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1932_  (.CLK(clknet_leaf_40_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0043_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0745_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1933_  (.CLK(clknet_3_6_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0044_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0746_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1934_  (.CLK(clknet_leaf_26_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0045_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0747_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1935_  (.CLK(clknet_leaf_32_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0046_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0748_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1936_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0047_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0749_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1937_  (.CLK(clknet_leaf_30_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0048_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0750_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1938_  (.CLK(clknet_leaf_40_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0049_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0751_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1939_  (.CLK(clknet_leaf_26_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0050_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0752_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1940_  (.CLK(clknet_leaf_25_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0051_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0753_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1941_  (.CLK(clknet_leaf_27_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0052_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0754_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1942_  (.CLK(clknet_leaf_22_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0053_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0755_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1943_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0054_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0756_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1944_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0055_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0757_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1945_  (.CLK(clknet_leaf_22_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0056_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0758_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1946_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0057_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0759_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1947_  (.CLK(clknet_leaf_22_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0058_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0760_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1948_  (.CLK(clknet_leaf_28_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0059_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0761_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1949_  (.CLK(clknet_leaf_28_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0060_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0762_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1950_  (.CLK(clknet_leaf_28_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0061_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0763_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1951_  (.CLK(clknet_leaf_28_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0062_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0764_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1952_  (.CLK(clknet_leaf_28_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0063_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0765_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1953_  (.CLK(clknet_leaf_27_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0064_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0766_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1954_  (.CLK(clknet_leaf_27_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0065_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0767_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1955_  (.CLK(clknet_leaf_27_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0066_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0768_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1956_  (.CLK(clknet_leaf_32_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0067_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0769_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1957_  (.CLK(clknet_3_6_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0068_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0770_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1958_  (.CLK(clknet_leaf_32_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0069_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0771_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1959_  (.CLK(clknet_leaf_32_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0070_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0772_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1960_  (.CLK(clknet_leaf_34_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0071_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0773_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1961_  (.CLK(clknet_leaf_34_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0072_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0774_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1962_  (.CLK(clknet_leaf_34_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0073_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0775_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1963_  (.CLK(clknet_leaf_39_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0074_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0776_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1964_  (.CLK(clknet_leaf_39_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0075_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0777_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1965_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0076_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0778_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1966_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0077_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0779_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1967_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0078_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0780_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1968_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0079_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0781_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1969_  (.CLK(clknet_leaf_35_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0080_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0782_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1970_  (.CLK(clknet_leaf_30_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0081_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0783_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1971_  (.CLK(clknet_leaf_30_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0082_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0784_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1972_  (.CLK(clknet_leaf_31_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0083_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0785_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1973_  (.CLK(clknet_leaf_29_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0084_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0786_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_rx._1974_  (.CLK(clknet_leaf_29_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_rx._0085_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_rx._0787_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1975_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net182),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1976_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1977_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1978_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1979_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1980_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1981_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1982_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0786_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1983_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net182),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1984_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1985_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1986_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1987_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1988_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1989_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1990_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0787_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1991_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1992_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net170),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1993_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1994_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1995_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net145),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1996_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net138),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1997_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net129),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1998_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0784_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._1999_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2000_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2001_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2002_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2003_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2004_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2005_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2006_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0785_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2007_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2008_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2009_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2010_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2011_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2012_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2013_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2014_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0758_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2015_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2016_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2017_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2018_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2019_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2020_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2021_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2022_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0760_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2023_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net180),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2024_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2025_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2026_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2027_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2028_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2029_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net131),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2030_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0754_ ),
    .D(net125),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2031_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2032_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net173),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2033_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2034_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2035_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2036_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net141),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2037_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2038_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0755_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2039_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net176),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2040_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net174),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2041_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2042_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2043_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net146),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2044_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2045_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2046_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0756_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2047_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2048_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2049_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net163),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2050_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net155),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2051_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net148),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2052_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2053_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2054_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0757_ ),
    .D(net122),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2055_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net177),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2056_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net167),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2057_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net160),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2058_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net152),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2059_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net144),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2060_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net135),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2061_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net128),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2062_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0759_ ),
    .D(net120),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2063_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net179),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2064_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2065_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net162),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2066_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net154),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2067_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net147),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2068_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2069_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net130),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2070_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0753_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2071_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2072_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2073_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2074_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2075_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2076_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2077_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2078_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0762_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2079_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net181),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2080_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net172),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2081_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net166),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2082_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net158),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2083_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2084_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net140),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2085_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net133),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2086_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0761_ ),
    .D(net124),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2087_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2088_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2089_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2090_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2091_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2092_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2093_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2094_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0724_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2095_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2096_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net171),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2097_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net165),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2098_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net157),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2099_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net150),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2100_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net139),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2101_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2102_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0722_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2103_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net178),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2104_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net174),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2105_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net164),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2106_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net156),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2107_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net149),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2108_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net142),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2109_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net132),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_rx._2110_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0723_ ),
    .D(net123),
    .Q(\u_usb_host.u_core.u_fifo_rx.ram[62][7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2111_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0013_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2112_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0014_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2113_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0015_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_rx._2114_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0016_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._2115_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0017_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_rx._2116_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_rx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_rx._0018_ ),
    .RESET_B(net401),
    .Q(\u_usb_host.u_core.u_fifo_rx.wr_ptr[5] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_tx._0788_  (.A(\u_usb_host.u_core.u_fifo_tx.count[6] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0443_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_tx._0789_  (.A(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0444_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_tx._0790_  (.A(\u_usb_host.u_core.u_fifo_tx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0445_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_tx._0791_  (.A(\u_usb_host.u_core.u_fifo_tx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_tx._0445_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0446_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_core.u_fifo_tx._0793_  (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0447_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_core.u_fifo_tx._0794_  (.A1(\u_usb_host.u_core.u_fifo_tx._0443_ ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0446_ ),
    .B1(net575),
    .X(\u_usb_host.u_core.u_fifo_tx._0448_ ));
 sky130_fd_sc_hd__o21ai_4 \u_usb_host.u_core.u_fifo_tx._0795_  (.A1(\u_usb_host.u_core.u_fifo_tx._0443_ ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0446_ ),
    .B1(net575),
    .Y(\u_usb_host.u_core.u_fifo_tx._0449_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_tx._0796_  (.A(net373),
    .B(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0450_ ));
 sky130_fd_sc_hd__and4_2 \u_usb_host.u_core.u_fifo_tx._0797_  (.A(net373),
    .B(net428),
    .C(net426),
    .D(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0451_ ));
 sky130_fd_sc_hd__nand3b_4 \u_usb_host.u_core.u_fifo_tx._0798_  (.A_N(net429),
    .B(net432),
    .C(\u_usb_host.u_core.u_fifo_tx._0451_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0452_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0799_  (.A(\u_usb_host.u_core.u_fifo_tx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0452_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0039_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0800_  (.A(net429),
    .B(net431),
    .X(\u_usb_host.u_core.u_fifo_tx._0453_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_core.u_fifo_tx._0801_  (.A(net428),
    .B(net426),
    .C(\u_usb_host.u_core.u_fifo_tx._0453_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0454_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_tx._0802_  (.A_N(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0455_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0803_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0455_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0456_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0804_  (.A(\u_usb_host.u_core.u_fifo_tx._0454_ ),
    .B(net104),
    .Y(\u_usb_host.u_core.u_fifo_tx._0042_ ));
 sky130_fd_sc_hd__nand4b_4 \u_usb_host.u_core.u_fifo_tx._0805_  (.A_N(net428),
    .B(net426),
    .C(net430),
    .D(net432),
    .Y(\u_usb_host.u_core.u_fifo_tx._0457_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0806_  (.A(\u_usb_host.u_core.u_fifo_tx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0458_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0807_  (.A(\u_usb_host.u_core.u_fifo_tx._0457_ ),
    .B(net103),
    .Y(\u_usb_host.u_core.u_fifo_tx._0037_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0808_  (.A(net429),
    .B(net431),
    .Y(\u_usb_host.u_core.u_fifo_tx._0459_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0809_  (.A(net429),
    .B(net431),
    .C(net428),
    .X(\u_usb_host.u_core.u_fifo_tx._0460_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_tx._0810_  (.A(net426),
    .B(\u_usb_host.u_core.u_fifo_tx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0461_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0811_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0041_ ));
 sky130_fd_sc_hd__or4b_2 \u_usb_host.u_core.u_fifo_tx._0812_  (.A(net431),
    .B(net428),
    .C(net426),
    .D_N(net429),
    .X(\u_usb_host.u_core.u_fifo_tx._0462_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0813_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0044_ ));
 sky130_fd_sc_hd__or4b_4 \u_usb_host.u_core.u_fifo_tx._0814_  (.A(net430),
    .B(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ),
    .C(net427),
    .D_N(net431),
    .X(\u_usb_host.u_core.u_fifo_tx._0463_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0815_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0043_ ));
 sky130_fd_sc_hd__or4bb_2 \u_usb_host.u_core.u_fifo_tx._0816_  (.A(net428),
    .B(net427),
    .C_N(net429),
    .D_N(net431),
    .X(\u_usb_host.u_core.u_fifo_tx._0464_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0817_  (.A(\u_usb_host.u_core.u_fifo_tx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0045_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_core.u_fifo_tx._0818_  (.A(net429),
    .B(net432),
    .C_N(\u_usb_host.u_core.u_fifo_tx._0451_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0465_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0819_  (.A(\u_usb_host.u_core.u_fifo_tx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0054_ ));
 sky130_fd_sc_hd__or4bb_2 \u_usb_host.u_core.u_fifo_tx._0820_  (.A(net432),
    .B(net427),
    .C_N(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ),
    .D_N(net430),
    .X(\u_usb_host.u_core.u_fifo_tx._0466_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0821_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0048_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0822_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0457_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0053_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_tx._0823_  (.A(net430),
    .B(net427),
    .C_N(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ),
    .D_N(net432),
    .X(\u_usb_host.u_core.u_fifo_tx._0467_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0824_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0047_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_tx._0825_  (.A(net431),
    .B(net428),
    .C_N(net426),
    .D_N(net429),
    .X(\u_usb_host.u_core.u_fifo_tx._0468_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0826_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0052_ ));
 sky130_fd_sc_hd__or4bb_4 \u_usb_host.u_core.u_fifo_tx._0827_  (.A(net429),
    .B(net428),
    .C_N(net426),
    .D_N(net431),
    .X(\u_usb_host.u_core.u_fifo_tx._0469_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0828_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0051_ ));
 sky130_fd_sc_hd__or3b_2 \u_usb_host.u_core.u_fifo_tx._0829_  (.A(\u_usb_host.u_core.u_fifo_tx._0453_ ),
    .B(net428),
    .C_N(net427),
    .X(\u_usb_host.u_core.u_fifo_tx._0470_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0830_  (.A(\u_usb_host.u_core.u_fifo_tx._0456_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0050_ ));
 sky130_fd_sc_hd__or4b_2 \u_usb_host.u_core.u_fifo_tx._0831_  (.A(net427),
    .B(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0453_ ),
    .D_N(net428),
    .X(\u_usb_host.u_core.u_fifo_tx._0471_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0832_  (.A(\u_usb_host.u_core.u_fifo_tx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0046_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_tx._0833_  (.A_N(net426),
    .B(\u_usb_host.u_core.u_fifo_tx._0460_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0472_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0834_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0049_ ));
 sky130_fd_sc_hd__nand3b_4 \u_usb_host.u_core.u_fifo_tx._0835_  (.A_N(net432),
    .B(\u_usb_host.u_core.u_fifo_tx._0451_ ),
    .C(net429),
    .Y(\u_usb_host.u_core.u_fifo_tx._0473_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0836_  (.A(\u_usb_host.u_core.u_fifo_tx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0040_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0837_  (.A(\u_usb_host.u_core.u_fifo_tx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0465_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0038_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0838_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0468_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0036_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0839_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0469_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0035_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0840_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0470_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0034_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0841_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0472_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0033_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_fifo_tx._0842_  (.A_N(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0474_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0843_  (.A(\u_usb_host.u_core.u_fifo_tx._0471_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0062_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core.u_fifo_tx._0844_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0464_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0061_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0845_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0475_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0846_  (.A(\u_usb_host.u_core.u_fifo_tx._0462_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0060_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0847_  (.A(\u_usb_host.u_core.u_fifo_tx._0463_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0475_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0059_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0848_  (.A(\u_usb_host.u_core.u_fifo_tx._0454_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0058_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0849_  (.A(net104),
    .B(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0057_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0850_  (.A(\u_usb_host.u_core.u_fifo_tx._0455_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0473_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0056_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0851_  (.A(\u_usb_host.u_core.u_fifo_tx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0455_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0055_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0852_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0466_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0032_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0853_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0467_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0031_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0854_  (.A(\u_usb_host.u_core.u_fifo_tx._0447_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0471_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0030_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0855_  (.A(net103),
    .B(\u_usb_host.u_core.u_fifo_tx._0464_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0029_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0856_  (.A(\u_usb_host.u_core.u_fifo_tx._0458_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0462_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0028_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0857_  (.A(\u_usb_host.u_core.u_fifo_tx._0458_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0463_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0027_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0858_  (.A(\u_usb_host.u_core.u_fifo_tx._0454_ ),
    .B(net103),
    .Y(\u_usb_host.u_core.u_fifo_tx._0026_ ));
 sky130_fd_sc_hd__o21a_2 \u_usb_host.u_core.u_fifo_tx._0860_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0446_ ),
    .B1(\u_usb_host.u_core.fifo_tx_pop_w ),
    .X(\u_usb_host.u_core.u_fifo_tx._0476_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_fifo_tx._0861_  (.A(\u_usb_host.u_core.u_fifo_tx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0477_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0862_  (.A(\u_usb_host.u_core.u_fifo_tx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0478_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_tx._0863_  (.A(\u_usb_host.u_core.u_fifo_tx.flush_i ),
    .B(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0025_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0864_  (.A(\u_usb_host.u_core.u_fifo_tx.flush_i ),
    .B(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0024_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0865_  (.A(\u_usb_host.u_core.u_fifo_tx.flush_i ),
    .B(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0023_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_tx._0866_  (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0479_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0867_  (.A(\u_usb_host.u_core.u_fifo_tx._0465_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0022_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0868_  (.A(\u_usb_host.u_core.u_fifo_tx._0473_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0021_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0869_  (.A(\u_usb_host.u_core.u_fifo_tx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0020_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0870_  (.A(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0480_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0871_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0480_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0019_ ));
 sky130_fd_sc_hd__or2_4 \u_usb_host.u_core.u_fifo_tx._0872_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0481_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0873_  (.A(\u_usb_host.u_core.u_fifo_tx._0462_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0076_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core.u_fifo_tx._0874_  (.A(\u_usb_host.u_core.u_fifo_tx._0450_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0463_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0075_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0875_  (.A(\u_usb_host.u_core.u_fifo_tx._0454_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0074_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0876_  (.A(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0073_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0877_  (.A(\u_usb_host.u_core.u_fifo_tx._0473_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0072_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0878_  (.A(\u_usb_host.u_core.u_fifo_tx._0452_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0071_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0879_  (.A(\u_usb_host.u_core.u_fifo_tx._0465_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0474_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0070_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0880_  (.A(\u_usb_host.u_core.u_fifo_tx._0457_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0069_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0881_  (.A(\u_usb_host.u_core.u_fifo_tx._0468_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0068_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0882_  (.A(\u_usb_host.u_core.u_fifo_tx._0469_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0067_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0883_  (.A(\u_usb_host.u_core.u_fifo_tx._0470_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0066_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0884_  (.A(\u_usb_host.u_core.u_fifo_tx._0466_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0064_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0885_  (.A(\u_usb_host.u_core.u_fifo_tx._0472_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0065_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0886_  (.A(\u_usb_host.u_core.u_fifo_tx._0467_ ),
    .B(net102),
    .Y(\u_usb_host.u_core.u_fifo_tx._0063_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0887_  (.A(\u_usb_host.u_core.u_fifo_tx._0472_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0081_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0888_  (.A(\u_usb_host.u_core.u_fifo_tx._0471_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0479_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0078_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0889_  (.A(\u_usb_host.u_core.u_fifo_tx._0466_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0080_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0890_  (.A(\u_usb_host.u_core.u_fifo_tx._0467_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0079_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0891_  (.A(\u_usb_host.u_core.u_fifo_tx._0464_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0077_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0892_  (.A(\u_usb_host.u_core.u_fifo_tx._0468_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0084_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0893_  (.A(\u_usb_host.u_core.u_fifo_tx._0457_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0085_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0894_  (.A(\u_usb_host.u_core.u_fifo_tx._0470_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0082_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0895_  (.A(\u_usb_host.u_core.u_fifo_tx._0469_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0481_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0083_ ));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_core.u_fifo_tx._0896_  (.A1(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B1_N(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0000_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_tx._0897_  (.A(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0482_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_fifo_tx._0898_  (.A0(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .A1(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .S(\u_usb_host.u_core.u_fifo_tx._0482_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0001_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_tx._0899_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0483_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0900_  (.A(\u_usb_host.u_core.u_fifo_tx._0444_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0483_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0484_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_tx._0901_  (.A(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .C(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0485_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_tx._0902_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0486_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._0903_  (.A1(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0485_ ),
    .A3(\u_usb_host.u_core.u_fifo_tx._0486_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0484_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0002_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0904_  (.A(\u_usb_host.u_core.u_fifo_tx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0444_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0487_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0905_  (.A(\u_usb_host.u_core.u_fifo_tx._0445_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0487_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0488_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_tx._0906_  (.A(\u_usb_host.u_core.u_fifo_tx.count[3] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .C(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .D(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0489_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_fifo_tx._0907_  (.A(\u_usb_host.u_core.u_fifo_tx._0489_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0490_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._0908_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx.count[0] ),
    .A3(\u_usb_host.u_core.u_fifo_tx.count[1] ),
    .B1(\u_usb_host.u_core.u_fifo_tx.count[3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0491_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._0909_  (.A1(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0490_ ),
    .A3(\u_usb_host.u_core.u_fifo_tx._0491_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0488_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0003_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_tx._0910_  (.A(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0445_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0492_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_tx._0911_  (.A(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0489_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0493_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_tx._0912_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0489_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0494_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_tx._0913_  (.A1_N(\u_usb_host.u_core.u_fifo_tx._0493_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_tx._0494_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0492_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0004_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_tx._0914_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0445_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx.count[5] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0495_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0915_  (.A(\u_usb_host.u_core.u_fifo_tx._0446_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0495_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0496_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0916_  (.A(\u_usb_host.u_core.u_fifo_tx.count[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.count[4] ),
    .C(\u_usb_host.u_core.u_fifo_tx._0489_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0497_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_tx._0917_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0493_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0498_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_fifo_tx._0918_  (.A1_N(\u_usb_host.u_core.u_fifo_tx._0497_ ),
    .A2_N(\u_usb_host.u_core.u_fifo_tx._0498_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0496_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0005_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_fifo_tx._0919_  (.A(\u_usb_host.u_core.u_fifo_tx._0443_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0497_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0499_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._0920_  (.A1(\u_usb_host.u_core.u_fifo_tx.count[6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0446_ ),
    .A3(\u_usb_host.u_core.u_fifo_tx._0478_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0499_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0477_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0006_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_tx._0921_  (.A_N(net440),
    .B(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0007_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0922_  (.A(net440),
    .B(net438),
    .Y(\u_usb_host.u_core.u_fifo_tx._0500_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0923_  (.A(net440),
    .B(net438),
    .X(\u_usb_host.u_core.u_fifo_tx._0501_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0924_  (.A(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0500_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0501_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0008_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_tx._0925_  (.A1(net440),
    .A2(net438),
    .B1(net436),
    .X(\u_usb_host.u_core.u_fifo_tx._0502_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_fifo_tx._0926_  (.A(net440),
    .B(net438),
    .C(net436),
    .Y(\u_usb_host.u_core.u_fifo_tx._0503_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0927_  (.A(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0502_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0503_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0009_ ));
 sky130_fd_sc_hd__and4b_2 \u_usb_host.u_core.u_fifo_tx._0928_  (.A_N(net433),
    .B(net435),
    .C(net437),
    .D(net439),
    .X(\u_usb_host.u_core.u_fifo_tx._0504_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_tx._0929_  (.A(net434),
    .B(\u_usb_host.u_core.u_fifo_tx._0503_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0505_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_fifo_tx._0930_  (.A1(net274),
    .A2(\u_usb_host.u_core.u_fifo_tx._0505_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0010_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_core.u_fifo_tx._0931_  (.A(net439),
    .B(net437),
    .C(net436),
    .D(net434),
    .X(\u_usb_host.u_core.u_fifo_tx._0506_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_fifo_tx._0932_  (.A1(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .A2(net272),
    .B1(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0507_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_fifo_tx._0933_  (.A1(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .A2(net272),
    .B1(\u_usb_host.u_core.u_fifo_tx._0507_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0011_ ));
 sky130_fd_sc_hd__and2b_2 \u_usb_host.u_core.u_fifo_tx._0934_  (.A_N(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ),
    .B(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0508_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_fifo_tx._0935_  (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0509_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_fifo_tx._0936_  (.A(net272),
    .B(net256),
    .Y(\u_usb_host.u_core.u_fifo_tx._0510_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_tx._0937_  (.A1(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .A2(net272),
    .B1(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0511_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0938_  (.A(\u_usb_host.u_core.u_fifo_tx._0476_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0510_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0511_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0012_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0939_  (.A(net431),
    .B(\u_usb_host.u_core.u_fifo_tx._0449_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0013_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0940_  (.A(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0453_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0459_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0014_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_fifo_tx._0941_  (.A1(net430),
    .A2(net431),
    .B1(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0512_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_core.u_fifo_tx._0942_  (.A_N(\u_usb_host.u_core.u_fifo_tx._0460_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0512_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0015_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_fifo_tx._0943_  (.A(net426),
    .B(\u_usb_host.u_core.u_fifo_tx._0460_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0513_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0944_  (.A(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0513_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0016_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_fifo_tx._0945_  (.A(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0461_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0514_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0946_  (.A(\u_usb_host.u_core.u_fifo_tx._0449_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0514_ ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0017_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._0947_  (.A1(net426),
    .A2(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ),
    .A3(\u_usb_host.u_core.u_fifo_tx._0460_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0515_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0948_  (.A(\u_usb_host.u_core.u_fifo_tx._0448_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0480_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0515_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0018_ ));
 sky130_fd_sc_hd__nor4_4 \u_usb_host.u_core.u_fifo_tx._0949_  (.A(net440),
    .B(net438),
    .C(net435),
    .D(net433),
    .Y(\u_usb_host.u_core.u_fifo_tx._0516_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_fifo_tx._0950_  (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ),
    .Y(\u_usb_host.u_core.u_fifo_tx._0517_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0951_  (.A(net243),
    .B(net239),
    .X(\u_usb_host.u_core.u_fifo_tx._0518_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_fifo_tx._0952_  (.A(net243),
    .B(net237),
    .Y(\u_usb_host.u_core.u_fifo_tx._0519_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_tx._0953_  (.A_N(net437),
    .B_N(net435),
    .C(net433),
    .D(net439),
    .X(\u_usb_host.u_core.u_fifo_tx._0520_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0954_  (.A(net268),
    .B(net232),
    .X(\u_usb_host.u_core.u_fifo_tx._0521_ ));
 sky130_fd_sc_hd__nor4b_1 \u_usb_host.u_core.u_fifo_tx._0955_  (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[0] ),
    .B(net436),
    .C(net434),
    .D_N(net437),
    .Y(\u_usb_host.u_core.u_fifo_tx._0522_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_fifo_tx._0956_  (.A_N(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ),
    .B(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0523_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0957_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][0] ),
    .B(net229),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_tx._0524_ ));
 sky130_fd_sc_hd__nor4b_4 \u_usb_host.u_core.u_fifo_tx._0958_  (.A(net440),
    .B(net438),
    .C(net435),
    .D_N(net433),
    .Y(\u_usb_host.u_core.u_fifo_tx._0525_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0959_  (.A(net268),
    .B(\u_usb_host.u_core.u_fifo_tx._0525_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0526_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_tx._0960_  (.A_N(net439),
    .B_N(net435),
    .C(net433),
    .D(net437),
    .X(\u_usb_host.u_core.u_fifo_tx._0527_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0961_  (.A(net237),
    .B(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0528_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_tx._0962_  (.A_N(net436),
    .B(net434),
    .C(net439),
    .D(net437),
    .X(\u_usb_host.u_core.u_fifo_tx._0529_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0963_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][0] ),
    .B(net218),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0530_ ));
 sky130_fd_sc_hd__nor4b_1 \u_usb_host.u_core.u_fifo_tx._0964_  (.A(net437),
    .B(net435),
    .C(net433),
    .D_N(net439),
    .Y(\u_usb_host.u_core.u_fifo_tx._0531_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0965_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][0] ),
    .B(net262),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0532_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0966_  (.A(net268),
    .B(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0533_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0967_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][0] ),
    .B(net251),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0534_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0968_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][0] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0535_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0969_  (.A(net237),
    .B(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0536_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0970_  (.A(net249),
    .B(\u_usb_host.u_core.u_fifo_tx._0525_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0537_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0971_  (.A(net237),
    .B(net232),
    .X(\u_usb_host.u_core.u_fifo_tx._0538_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0972_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][0] ),
    .B(net264),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0539_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0973_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][0] ),
    .B(net255),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0540_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0974_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][0] ),
    .B(net232),
    .C(net218),
    .X(\u_usb_host.u_core.u_fifo_tx._0541_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0975_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][0] ),
    .B(net263),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0542_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0976_  (.A(net239),
    .B(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0543_ ));
 sky130_fd_sc_hd__and4bb_2 \u_usb_host.u_core.u_fifo_tx._0977_  (.A_N(net435),
    .B_N(net433),
    .C(net439),
    .D(net437),
    .X(\u_usb_host.u_core.u_fifo_tx._0544_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0978_  (.A(net239),
    .B(\u_usb_host.u_core.u_fifo_tx._0544_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0545_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0979_  (.A(net268),
    .B(\u_usb_host.u_core.u_fifo_tx._0544_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0546_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0980_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][0] ),
    .B(net243),
    .C(net219),
    .X(\u_usb_host.u_core.u_fifo_tx._0547_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0981_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][0] ),
    .B(net222),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0548_ ));
 sky130_fd_sc_hd__nor4b_1 \u_usb_host.u_core.u_fifo_tx._0982_  (.A(\u_usb_host.u_core.u_fifo_tx.rd_ptr[0] ),
    .B(net437),
    .C(net434),
    .D_N(net436),
    .Y(\u_usb_host.u_core.u_fifo_tx._0549_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0983_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][0] ),
    .B(net247),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0550_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0984_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][0] ),
    .B(net244),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0551_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0985_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][0] ),
    .B(net257),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0552_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0986_  (.A(net239),
    .B(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0553_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0987_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][0] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0554_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0988_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][0] ),
    .B(net239),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0555_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0989_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][0] ),
    .B(net248),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0556_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0990_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][0] ),
    .B(net220),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0557_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0991_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][0] ),
    .B(net225),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0558_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0992_  (.A(net268),
    .B(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0559_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0993_  (.A(net218),
    .B(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0560_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._0994_  (.A(net274),
    .B(net268),
    .X(\u_usb_host.u_core.u_fifo_tx._0561_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0995_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][0] ),
    .B(net272),
    .C(net254),
    .X(\u_usb_host.u_core.u_fifo_tx._0562_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_tx._0996_  (.A_N(net440),
    .B_N(net438),
    .C(net435),
    .D(net433),
    .X(\u_usb_host.u_core.u_fifo_tx._0563_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0997_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][0] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0564_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._0998_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][0] ),
    .B(net220),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0565_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_tx._0999_  (.A_N(net438),
    .B(net436),
    .C(net434),
    .D(net439),
    .X(\u_usb_host.u_core.u_fifo_tx._0566_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1000_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][0] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0567_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1001_  (.A(net274),
    .B(net250),
    .X(\u_usb_host.u_core.u_fifo_tx._0568_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1002_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][0] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0569_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1003_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][0] ),
    .B(net270),
    .C(net265),
    .X(\u_usb_host.u_core.u_fifo_tx._0570_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_tx._1004_  (.A_N(\u_usb_host.u_core.u_fifo_tx.rd_ptr[1] ),
    .B_N(net434),
    .C(net436),
    .D(net439),
    .X(\u_usb_host.u_core.u_fifo_tx._0571_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1005_  (.A(net237),
    .B(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0572_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_fifo_tx._1006_  (.A_N(net440),
    .B(net438),
    .C(net435),
    .D(net433),
    .X(\u_usb_host.u_core.u_fifo_tx._0573_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1007_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][0] ),
    .B(net271),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0574_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_fifo_tx._1008_  (.A_N(net439),
    .B_N(net433),
    .C(net435),
    .D(net437),
    .X(\u_usb_host.u_core.u_fifo_tx._0575_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1009_  (.A(net238),
    .B(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0576_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1010_  (.A(net237),
    .B(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0577_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1011_  (.A(net274),
    .B(net239),
    .X(\u_usb_host.u_core.u_fifo_tx._0578_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1012_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][0] ),
    .B(net251),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0579_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1013_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][0] ),
    .B(net214),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0580_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1014_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][0] ),
    .B(net274),
    .C(net225),
    .X(\u_usb_host.u_core.u_fifo_tx._0581_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1015_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][0] ),
    .B(net267),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0582_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1016_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][0] ),
    .B(net252),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0583_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1017_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][0] ),
    .B(net225),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0584_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1018_  (.A(net250),
    .B(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0585_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1019_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][0] ),
    .B(net267),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0586_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1020_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][0] ),
    .B(net247),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0587_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1021_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][0] ),
    .B(net234),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0588_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1022_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][0] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0589_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1023_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][0] ),
    .B(net255),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0590_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_fifo_tx._1024_  (.A(net267),
    .B(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0591_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1025_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][0] ),
    .B(net226),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0592_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1026_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0593_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1027_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[14][0] ),
    .A2(net234),
    .A3(net185),
    .B1(\u_usb_host.u_core.u_fifo_tx._0588_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0535_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0594_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1028_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0595_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1029_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0596_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1030_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][0] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0595_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0597_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1031_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][0] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0596_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0598_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1032_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][0] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0593_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0599_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1033_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][0] ),
    .A2(net260),
    .A3(net192),
    .B1(\u_usb_host.u_core.u_fifo_tx._0589_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0600_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1034_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][0] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0600_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0547_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0601_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1035_  (.A(\u_usb_host.u_core.u_fifo_tx._0597_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0598_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0599_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0601_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0602_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_tx._1036_  (.A(\u_usb_host.u_core.u_fifo_tx._0551_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0567_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0569_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0580_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0603_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1037_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0564_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0530_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0541_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0604_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1038_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0542_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0539_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0532_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0605_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1039_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0586_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0582_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0570_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0606_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1040_  (.A(\u_usb_host.u_core.u_fifo_tx._0603_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0604_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0605_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0606_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0607_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1041_  (.A(\u_usb_host.u_core.u_fifo_tx._0540_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0555_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0562_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0590_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0608_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1042_  (.A(\u_usb_host.u_core.u_fifo_tx._0534_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0552_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0579_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0583_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0609_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1043_  (.A(\u_usb_host.u_core.u_fifo_tx._0524_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0548_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0557_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0565_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0610_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1044_  (.A(\u_usb_host.u_core.u_fifo_tx._0558_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0581_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0584_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0592_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0611_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1045_  (.A(\u_usb_host.u_core.u_fifo_tx._0608_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0609_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0610_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0611_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0612_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1046_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0613_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1047_  (.A(\u_usb_host.u_core.u_fifo_tx._0550_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0554_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0556_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0587_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0614_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1048_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0613_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0614_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0615_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1049_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0616_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1050_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][0] ),
    .A2(net237),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][0] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0617_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1051_  (.A(\u_usb_host.u_core.u_fifo_tx._0574_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0594_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0616_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0617_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0618_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1052_  (.A(\u_usb_host.u_core.u_fifo_tx._0607_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0612_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0615_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0618_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0619_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1053_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][0] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0602_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0619_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[0] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1054_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][1] ),
    .B(net227),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0620_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1055_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][1] ),
    .B(net220),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0621_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1056_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][1] ),
    .B(net216),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0622_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1057_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][1] ),
    .B(net262),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0623_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1058_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][1] ),
    .B(net251),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0624_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1059_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][1] ),
    .B(net223),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0625_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1060_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][1] ),
    .B(net246),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0626_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1061_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][1] ),
    .B(net264),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0627_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1062_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][1] ),
    .B(net254),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0628_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1063_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][1] ),
    .B(net244),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0629_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1064_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][1] ),
    .B(net262),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0630_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1065_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][1] ),
    .B(net243),
    .C(net219),
    .X(\u_usb_host.u_core.u_fifo_tx._0631_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1066_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][1] ),
    .B(net252),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0632_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1067_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][1] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0633_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1068_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][1] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0634_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1069_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][1] ),
    .B(net239),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0635_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1070_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][1] ),
    .B(net232),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_tx._0636_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1071_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][1] ),
    .B(net230),
    .C(net222),
    .X(\u_usb_host.u_core.u_fifo_tx._0637_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1072_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][1] ),
    .B(net272),
    .C(net253),
    .X(\u_usb_host.u_core.u_fifo_tx._0638_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1073_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][1] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0639_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1074_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][1] ),
    .B(net253),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0640_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1075_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][1] ),
    .B(net267),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0641_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1076_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][1] ),
    .B(net225),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0642_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1077_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[14][1] ),
    .B(net235),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0643_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1078_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][1] ),
    .B(net269),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0644_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1079_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][1] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0645_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1080_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][1] ),
    .B(net250),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0646_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1081_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][1] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0647_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1082_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][1] ),
    .B(net270),
    .C(net266),
    .X(\u_usb_host.u_core.u_fifo_tx._0648_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1083_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][1] ),
    .B(net227),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0649_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1084_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][1] ),
    .B(net214),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0650_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1085_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][1] ),
    .B(net251),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0651_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1086_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][1] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0652_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1087_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][1] ),
    .B(net246),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0653_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1088_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][1] ),
    .B(net246),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0654_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1089_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][1] ),
    .B(net265),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0655_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1090_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][1] ),
    .B(net222),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0656_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1091_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][1] ),
    .B(net274),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_tx._0657_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1092_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0658_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1093_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[13][1] ),
    .A2(net235),
    .A3(net194),
    .B1(\u_usb_host.u_core.u_fifo_tx._0634_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0643_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0659_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1094_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0660_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1095_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0661_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1096_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][1] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0660_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0662_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1097_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][1] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0661_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0663_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1098_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][1] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0658_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0664_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1099_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][1] ),
    .A2(net260),
    .A3(net192),
    .B1(\u_usb_host.u_core.u_fifo_tx._0645_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0665_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1100_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][1] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0631_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0665_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0666_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1101_  (.A(\u_usb_host.u_core.u_fifo_tx._0662_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0663_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0664_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0666_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0667_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1102_  (.A(\u_usb_host.u_core.u_fifo_tx._0629_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0647_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0650_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0652_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0668_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1103_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0622_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0636_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0639_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0669_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1104_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0623_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0627_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0630_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0670_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1105_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0641_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0648_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0655_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0671_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1106_  (.A(\u_usb_host.u_core.u_fifo_tx._0668_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0669_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0670_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0671_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0672_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1107_  (.A(\u_usb_host.u_core.u_fifo_tx._0628_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0635_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0638_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0640_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0673_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1108_  (.A(\u_usb_host.u_core.u_fifo_tx._0624_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0632_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0646_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0651_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0674_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1109_  (.A(\u_usb_host.u_core.u_fifo_tx._0621_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0625_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0637_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0656_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0675_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1110_  (.A(\u_usb_host.u_core.u_fifo_tx._0620_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0642_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0649_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0657_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0676_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1111_  (.A(\u_usb_host.u_core.u_fifo_tx._0673_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0674_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0675_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0676_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0677_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1112_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0678_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1113_  (.A(\u_usb_host.u_core.u_fifo_tx._0626_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0633_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0653_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0654_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0679_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1114_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0678_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0679_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0680_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1115_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0681_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1116_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][1] ),
    .A2(net236),
    .A3(net196),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][1] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0682_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_tx._1117_  (.A(\u_usb_host.u_core.u_fifo_tx._0644_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0659_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0681_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0682_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0683_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1118_  (.A(\u_usb_host.u_core.u_fifo_tx._0672_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0677_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0680_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0683_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0684_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1119_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][1] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0667_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0684_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[1] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1120_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][2] ),
    .B(net230),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_tx._0685_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1121_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][2] ),
    .B(net217),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0686_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1122_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][2] ),
    .B(net262),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0687_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1123_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][2] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0688_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1124_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][2] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0689_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1125_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][2] ),
    .B(net264),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0690_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1126_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][2] ),
    .B(net255),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0691_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1127_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][2] ),
    .B(net232),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_tx._0692_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1128_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][2] ),
    .B(net262),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0693_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1129_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][2] ),
    .B(net243),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_tx._0694_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1130_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][2] ),
    .B(net252),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0695_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1131_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][2] ),
    .B(net246),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0696_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1132_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][2] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0697_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1133_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][2] ),
    .B(net251),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0698_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1134_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][2] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0699_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1135_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][2] ),
    .B(net239),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0700_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1136_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][2] ),
    .B(net246),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0701_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1137_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][2] ),
    .B(net220),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0702_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1138_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][2] ),
    .B(net227),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0703_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1139_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][2] ),
    .B(net272),
    .C(net254),
    .X(\u_usb_host.u_core.u_fifo_tx._0704_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1140_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][2] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0705_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1141_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][2] ),
    .B(net220),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0706_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1142_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][2] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0707_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1143_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][2] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0708_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1144_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][2] ),
    .B(net270),
    .C(net265),
    .X(\u_usb_host.u_core.u_fifo_tx._0709_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1145_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][2] ),
    .B(net269),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0710_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1146_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][2] ),
    .B(net250),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0711_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1147_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][2] ),
    .B(net213),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0712_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1148_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][2] ),
    .B(net274),
    .C(net227),
    .X(\u_usb_host.u_core.u_fifo_tx._0713_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1149_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][2] ),
    .B(net267),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0714_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1150_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][2] ),
    .B(net251),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0715_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1151_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][2] ),
    .B(net224),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0716_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1152_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][2] ),
    .B(net265),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0717_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1153_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][2] ),
    .B(net247),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0718_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1154_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][2] ),
    .B(net234),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0719_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1155_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][2] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0720_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1156_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][2] ),
    .B(net227),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0086_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1157_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][2] ),
    .B(net255),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0087_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1158_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0088_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1159_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[14][2] ),
    .A2(net234),
    .A3(net185),
    .B1(\u_usb_host.u_core.u_fifo_tx._0689_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0719_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0089_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1160_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0090_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1161_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0091_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1162_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][2] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0090_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0092_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1163_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][2] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0091_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0093_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1164_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][2] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0088_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0094_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1165_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][2] ),
    .A2(net260),
    .A3(net194),
    .B1(\u_usb_host.u_core.u_fifo_tx._0720_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0095_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1166_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][2] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0694_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0095_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0096_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1167_  (.A(\u_usb_host.u_core.u_fifo_tx._0092_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0093_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0094_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0096_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0097_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1168_  (.A(\u_usb_host.u_core.u_fifo_tx._0697_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0707_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0708_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0712_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0098_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1169_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0686_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0692_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0705_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0099_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1170_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0687_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0690_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0693_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0100_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1171_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0709_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0714_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0717_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0101_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1172_  (.A(\u_usb_host.u_core.u_fifo_tx._0098_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0099_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0100_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0101_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0102_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1173_  (.A(\u_usb_host.u_core.u_fifo_tx._0691_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0700_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0704_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0087_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0103_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1174_  (.A(\u_usb_host.u_core.u_fifo_tx._0695_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0698_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0711_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0715_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0104_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1175_  (.A(\u_usb_host.u_core.u_fifo_tx._0685_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0688_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0702_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0706_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0105_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1176_  (.A(\u_usb_host.u_core.u_fifo_tx._0703_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0713_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0716_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0086_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0106_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1177_  (.A(\u_usb_host.u_core.u_fifo_tx._0103_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0104_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0105_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0106_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0107_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1178_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0108_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1179_  (.A(\u_usb_host.u_core.u_fifo_tx._0696_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0699_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0701_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0718_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0109_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1180_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0108_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0109_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0110_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1181_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0111_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1182_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][2] ),
    .A2(net236),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][2] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0112_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1183_  (.A(\u_usb_host.u_core.u_fifo_tx._0710_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0089_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0111_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0112_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0113_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1184_  (.A(\u_usb_host.u_core.u_fifo_tx._0102_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0107_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0110_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0113_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0114_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1185_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][2] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0097_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0114_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[2] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1186_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][3] ),
    .B(net221),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0115_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1187_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][3] ),
    .B(net217),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0116_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1188_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][3] ),
    .B(net262),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0117_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1189_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][3] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0118_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1190_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][3] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0119_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1191_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][3] ),
    .B(net264),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0120_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1192_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][3] ),
    .B(net253),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0121_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1193_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][3] ),
    .B(net232),
    .C(net217),
    .X(\u_usb_host.u_core.u_fifo_tx._0122_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1194_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][3] ),
    .B(net262),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0123_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1195_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][3] ),
    .B(net243),
    .C(net219),
    .X(\u_usb_host.u_core.u_fifo_tx._0124_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1196_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][3] ),
    .B(net251),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0125_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1197_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][3] ),
    .B(net247),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0126_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1198_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][3] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0127_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1199_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][3] ),
    .B(net257),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0128_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1200_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][3] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0129_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1201_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][3] ),
    .B(net239),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0130_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1202_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][3] ),
    .B(net246),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0131_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1203_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][3] ),
    .B(net230),
    .C(net222),
    .X(\u_usb_host.u_core.u_fifo_tx._0132_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1204_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][3] ),
    .B(net224),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0133_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1205_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][3] ),
    .B(net272),
    .C(net254),
    .X(\u_usb_host.u_core.u_fifo_tx._0134_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1206_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][3] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0135_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1207_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][3] ),
    .B(net224),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0136_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1208_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][3] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0137_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1209_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][3] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0138_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1210_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][3] ),
    .B(net270),
    .C(net265),
    .X(\u_usb_host.u_core.u_fifo_tx._0139_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1211_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][3] ),
    .B(net271),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0140_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1212_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][3] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0141_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1213_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][3] ),
    .B(net251),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0142_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1214_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][3] ),
    .B(net213),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0143_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1215_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][3] ),
    .B(net253),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0144_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1216_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][3] ),
    .B(net267),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0145_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1217_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][3] ),
    .B(net251),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0146_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1218_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][3] ),
    .B(net224),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0147_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1219_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][3] ),
    .B(net265),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0148_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1220_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][3] ),
    .B(net222),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0149_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1221_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][3] ),
    .B(net247),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0150_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1222_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][3] ),
    .B(net234),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0151_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1223_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][3] ),
    .B(net274),
    .C(net224),
    .X(\u_usb_host.u_core.u_fifo_tx._0152_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1224_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0153_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1225_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[14][3] ),
    .A2(net234),
    .A3(net185),
    .B1(\u_usb_host.u_core.u_fifo_tx._0119_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0151_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0154_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1226_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0155_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1227_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0156_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1228_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][3] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0155_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0157_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1229_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][3] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0156_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0158_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1230_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][3] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0153_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0159_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1231_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][3] ),
    .A2(net260),
    .A3(net192),
    .B1(\u_usb_host.u_core.u_fifo_tx._0141_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0160_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1232_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][3] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0124_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0160_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0161_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1233_  (.A(\u_usb_host.u_core.u_fifo_tx._0157_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0158_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0159_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0161_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0162_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1234_  (.A(\u_usb_host.u_core.u_fifo_tx._0127_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0137_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0138_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0143_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0163_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1235_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0116_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0122_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0135_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0164_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1236_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0117_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0120_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0123_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0165_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1237_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0139_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0145_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0148_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0166_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1238_  (.A(\u_usb_host.u_core.u_fifo_tx._0163_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0164_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0165_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0166_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0167_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1239_  (.A(\u_usb_host.u_core.u_fifo_tx._0121_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0130_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0134_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0144_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0168_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1240_  (.A(\u_usb_host.u_core.u_fifo_tx._0125_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0128_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0142_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0146_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0169_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1241_  (.A(\u_usb_host.u_core.u_fifo_tx._0115_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0118_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0132_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0149_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0170_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1242_  (.A(\u_usb_host.u_core.u_fifo_tx._0133_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0136_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0147_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0152_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0171_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1243_  (.A(\u_usb_host.u_core.u_fifo_tx._0168_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0169_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0170_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0171_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0172_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1244_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0173_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1245_  (.A(\u_usb_host.u_core.u_fifo_tx._0126_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0129_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0131_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0150_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0174_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1246_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0173_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0174_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0175_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1247_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0176_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1248_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][3] ),
    .A2(net238),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][3] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0177_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1249_  (.A(\u_usb_host.u_core.u_fifo_tx._0140_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0154_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0176_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0177_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0178_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1250_  (.A(\u_usb_host.u_core.u_fifo_tx._0167_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0172_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0175_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0178_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0179_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1251_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][3] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0162_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0179_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[3] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1252_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][4] ),
    .B(net263),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0180_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1253_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][4] ),
    .B(net230),
    .C(net222),
    .X(\u_usb_host.u_core.u_fifo_tx._0181_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1254_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][4] ),
    .B(net257),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0182_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1255_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][4] ),
    .B(net217),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0183_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1256_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][4] ),
    .B(net240),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0184_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1257_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][4] ),
    .B(net225),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0185_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1258_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][4] ),
    .B(net247),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0186_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1259_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][4] ),
    .B(net263),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0187_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1260_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][4] ),
    .B(net253),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0188_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1261_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][4] ),
    .B(net243),
    .C(net213),
    .X(\u_usb_host.u_core.u_fifo_tx._0189_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1262_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][4] ),
    .B(net263),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0190_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1263_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][4] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0191_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1264_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][4] ),
    .B(net257),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0192_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1265_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][4] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0193_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1266_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][4] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0194_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1267_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][4] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0195_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1268_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][4] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0196_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1269_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][4] ),
    .B(net221),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0197_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1270_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][4] ),
    .B(net232),
    .C(net218),
    .X(\u_usb_host.u_core.u_fifo_tx._0198_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1271_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][4] ),
    .B(net222),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0199_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1272_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][4] ),
    .B(net272),
    .C(net253),
    .X(\u_usb_host.u_core.u_fifo_tx._0200_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1273_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][4] ),
    .B(net246),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0201_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1274_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[14][4] ),
    .B(net234),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0202_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1275_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][4] ),
    .B(net270),
    .C(net266),
    .X(\u_usb_host.u_core.u_fifo_tx._0203_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1276_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][4] ),
    .B(net235),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0204_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1277_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][4] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0205_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1278_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][4] ),
    .B(net269),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0206_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1279_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0207_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1280_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][4] ),
    .B(net268),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0208_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1281_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][4] ),
    .B(net249),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0209_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1282_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][4] ),
    .B(net214),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0210_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1283_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][4] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0211_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1284_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][4] ),
    .B(net225),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0212_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1285_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][4] ),
    .B(net274),
    .C(net226),
    .X(\u_usb_host.u_core.u_fifo_tx._0213_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1286_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][4] ),
    .B(net252),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0214_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1287_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][4] ),
    .B(net247),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0215_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1288_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][4] ),
    .B(net253),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0216_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1289_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][4] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0217_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1290_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][4] ),
    .B(net226),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0218_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1291_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][4] ),
    .B(net265),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0219_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1292_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0220_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1293_  (.A(\u_usb_host.u_core.u_fifo_tx._0195_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0202_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0204_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0206_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0221_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1294_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0222_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1295_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][4] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0207_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0223_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1296_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][4] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0222_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0224_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1297_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][4] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0220_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0225_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1298_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][4] ),
    .A2(net259),
    .A3(net193),
    .B1(\u_usb_host.u_core.u_fifo_tx._0217_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0226_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1299_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][4] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0189_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0226_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0227_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1300_  (.A(\u_usb_host.u_core.u_fifo_tx._0223_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0224_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0225_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0227_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0228_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1301_  (.A(\u_usb_host.u_core.u_fifo_tx._0193_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0196_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0210_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0211_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0229_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1302_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0183_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0198_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0205_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0230_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1303_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0180_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0187_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0190_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0231_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1304_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0203_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0208_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0219_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0232_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1305_  (.A(\u_usb_host.u_core.u_fifo_tx._0229_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0230_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0231_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0232_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0233_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1306_  (.A(\u_usb_host.u_core.u_fifo_tx._0184_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0188_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0200_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0216_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0234_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1307_  (.A(\u_usb_host.u_core.u_fifo_tx._0182_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0192_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0209_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0214_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0235_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1308_  (.A(\u_usb_host.u_core.u_fifo_tx._0181_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0191_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0197_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0199_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0236_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1309_  (.A(\u_usb_host.u_core.u_fifo_tx._0185_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0212_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0213_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0218_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0237_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1310_  (.A(\u_usb_host.u_core.u_fifo_tx._0234_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0235_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0236_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0237_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0238_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1311_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0239_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1312_  (.A(\u_usb_host.u_core.u_fifo_tx._0186_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0194_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0201_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0215_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0240_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1313_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0239_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0240_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0241_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1314_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0242_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1315_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][4] ),
    .A2(net237),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][4] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0243_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_tx._1316_  (.A(\u_usb_host.u_core.u_fifo_tx._0221_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0242_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0243_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0244_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1317_  (.A(\u_usb_host.u_core.u_fifo_tx._0233_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0238_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0241_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0244_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0245_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1318_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][4] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0228_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0245_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[4] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1319_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][5] ),
    .B(net230),
    .C(net220),
    .X(\u_usb_host.u_core.u_fifo_tx._0246_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1320_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][5] ),
    .B(net257),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0247_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1321_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][5] ),
    .B(net218),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0248_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1322_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][5] ),
    .B(net240),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0249_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1323_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][5] ),
    .B(net227),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0250_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1324_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][5] ),
    .B(net248),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0251_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1325_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][5] ),
    .B(net263),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0252_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1326_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][5] ),
    .B(net253),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0253_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1327_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][5] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0254_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1328_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][5] ),
    .B(net263),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0255_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1329_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][5] ),
    .B(net262),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0256_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1330_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][5] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0257_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1331_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][5] ),
    .B(net257),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0258_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1332_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][5] ),
    .B(net215),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0259_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1333_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][5] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0260_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1334_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][5] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0261_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1335_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][5] ),
    .B(net232),
    .C(net218),
    .X(\u_usb_host.u_core.u_fifo_tx._0262_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1336_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][5] ),
    .B(net221),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0263_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1337_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][5] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0516_ ),
    .C(net215),
    .X(\u_usb_host.u_core.u_fifo_tx._0264_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1338_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][5] ),
    .B(net222),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0265_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1339_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][5] ),
    .B(net273),
    .C(net253),
    .X(\u_usb_host.u_core.u_fifo_tx._0266_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1340_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][5] ),
    .B(net268),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0267_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1341_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][5] ),
    .B(net235),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0268_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1342_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][5] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0269_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1343_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[14][5] ),
    .B(net234),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0270_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1344_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][5] ),
    .B(net269),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0271_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1345_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0272_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1346_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][5] ),
    .B(net249),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0273_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1347_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][5] ),
    .B(net270),
    .C(net215),
    .X(\u_usb_host.u_core.u_fifo_tx._0274_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1348_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][5] ),
    .B(net271),
    .C(net266),
    .X(\u_usb_host.u_core.u_fifo_tx._0275_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1349_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][5] ),
    .B(net274),
    .C(net226),
    .X(\u_usb_host.u_core.u_fifo_tx._0276_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1350_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][5] ),
    .B(net252),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0277_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1351_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][5] ),
    .B(net215),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0278_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1352_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][5] ),
    .B(net225),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0279_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1353_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][5] ),
    .B(net247),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0280_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1354_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][5] ),
    .B(net256),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0281_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1355_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][5] ),
    .B(net246),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0282_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1356_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][5] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0283_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1357_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][5] ),
    .B(net226),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0284_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1358_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][5] ),
    .B(net267),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0285_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1359_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0286_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1360_  (.A(\u_usb_host.u_core.u_fifo_tx._0261_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0268_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0270_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0271_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0287_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1361_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0288_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1362_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][5] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0272_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0289_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1363_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][5] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0288_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0290_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1364_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][5] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0286_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0291_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1365_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][5] ),
    .A2(net260),
    .A3(net194),
    .B1(\u_usb_host.u_core.u_fifo_tx._0283_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0292_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1366_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][5] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0264_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0292_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0293_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1367_  (.A(\u_usb_host.u_core.u_fifo_tx._0289_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0290_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0291_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0293_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0294_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1368_  (.A(\u_usb_host.u_core.u_fifo_tx._0254_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0259_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0274_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0278_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0295_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1369_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0248_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0262_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0269_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0296_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1370_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0252_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0255_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0256_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0297_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1371_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0267_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0275_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0285_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0298_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1372_  (.A(\u_usb_host.u_core.u_fifo_tx._0295_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0296_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0297_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0298_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0299_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1373_  (.A(\u_usb_host.u_core.u_fifo_tx._0249_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0253_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0266_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0281_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0300_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1374_  (.A(\u_usb_host.u_core.u_fifo_tx._0247_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0258_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0273_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0277_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0301_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1375_  (.A(\u_usb_host.u_core.u_fifo_tx._0246_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0257_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0263_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0265_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0302_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1376_  (.A(\u_usb_host.u_core.u_fifo_tx._0250_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0276_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0279_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0284_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0303_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1377_  (.A(\u_usb_host.u_core.u_fifo_tx._0300_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0301_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0302_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0303_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0304_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1378_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0305_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1379_  (.A(\u_usb_host.u_core.u_fifo_tx._0251_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0260_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0280_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0282_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0306_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1380_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0305_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0306_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0307_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1381_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0308_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1382_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][5] ),
    .A2(net237),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][5] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0309_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_tx._1383_  (.A(\u_usb_host.u_core.u_fifo_tx._0287_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0308_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0309_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0310_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1384_  (.A(\u_usb_host.u_core.u_fifo_tx._0299_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0304_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0307_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0310_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0311_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1385_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][5] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0294_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0311_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[5] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1386_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][6] ),
    .B(net230),
    .C(net221),
    .X(\u_usb_host.u_core.u_fifo_tx._0312_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1387_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][6] ),
    .B(net257),
    .C(net210),
    .X(\u_usb_host.u_core.u_fifo_tx._0313_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1388_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][6] ),
    .B(net218),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0314_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1389_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][6] ),
    .B(net257),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0315_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1390_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][6] ),
    .B(net225),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0316_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1391_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][6] ),
    .B(net248),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0317_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1392_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][6] ),
    .B(net263),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0318_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1393_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][6] ),
    .B(net255),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0319_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1394_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][6] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0320_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1395_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][6] ),
    .B(net263),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0321_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1396_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][6] ),
    .B(net263),
    .C(net206),
    .X(\u_usb_host.u_core.u_fifo_tx._0322_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1397_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][6] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0323_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1398_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][6] ),
    .B(net240),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0324_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1399_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][6] ),
    .B(net215),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0325_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1400_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][6] ),
    .B(net248),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0326_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1401_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][6] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0327_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1402_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][6] ),
    .B(net232),
    .C(net218),
    .X(\u_usb_host.u_core.u_fifo_tx._0328_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1403_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][6] ),
    .B(net221),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0329_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1404_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][6] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0516_ ),
    .C(net215),
    .X(\u_usb_host.u_core.u_fifo_tx._0330_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1405_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][6] ),
    .B(net220),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0331_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1406_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][6] ),
    .B(net273),
    .C(net254),
    .X(\u_usb_host.u_core.u_fifo_tx._0332_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1407_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][6] ),
    .B(net267),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0333_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1408_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[13][6] ),
    .B(net235),
    .C(net192),
    .X(\u_usb_host.u_core.u_fifo_tx._0334_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1409_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][6] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0335_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1410_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[14][6] ),
    .B(net234),
    .C(net185),
    .X(\u_usb_host.u_core.u_fifo_tx._0336_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1411_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][6] ),
    .B(net270),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0337_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1412_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0338_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1413_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][6] ),
    .B(net258),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0339_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1414_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][6] ),
    .B(net270),
    .C(net215),
    .X(\u_usb_host.u_core.u_fifo_tx._0340_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1415_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][6] ),
    .B(net271),
    .C(net265),
    .X(\u_usb_host.u_core.u_fifo_tx._0341_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1416_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][6] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0504_ ),
    .C(net225),
    .X(\u_usb_host.u_core.u_fifo_tx._0342_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1417_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][6] ),
    .B(net251),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0343_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1418_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][6] ),
    .B(net215),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0344_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1419_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][6] ),
    .B(net225),
    .C(net184),
    .X(\u_usb_host.u_core.u_fifo_tx._0345_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1420_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][6] ),
    .B(net247),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0346_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1421_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][6] ),
    .B(net255),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0347_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1422_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][6] ),
    .B(net246),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0348_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1423_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][6] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0349_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1424_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][6] ),
    .B(net226),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0350_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1425_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][6] ),
    .B(net267),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0351_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1426_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0352_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1427_  (.A(\u_usb_host.u_core.u_fifo_tx._0327_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0334_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0336_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0337_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0353_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1428_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0354_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1429_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][6] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0338_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0355_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1430_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][6] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0354_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0356_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1431_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][6] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0352_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0357_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1432_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][6] ),
    .A2(net259),
    .A3(net194),
    .B1(\u_usb_host.u_core.u_fifo_tx._0349_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0358_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1433_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][6] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0330_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0358_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0359_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1434_  (.A(\u_usb_host.u_core.u_fifo_tx._0355_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0356_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0357_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0359_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0360_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1435_  (.A(\u_usb_host.u_core.u_fifo_tx._0320_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0325_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0340_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0344_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0361_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1436_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0314_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0328_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0335_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0362_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1437_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0318_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0321_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0322_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0363_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1438_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0333_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0341_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0351_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0364_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1439_  (.A(\u_usb_host.u_core.u_fifo_tx._0361_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0362_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0363_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0364_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0365_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1440_  (.A(\u_usb_host.u_core.u_fifo_tx._0319_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0324_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0332_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0347_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0366_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1441_  (.A(\u_usb_host.u_core.u_fifo_tx._0313_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0315_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0339_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0343_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0367_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1442_  (.A(\u_usb_host.u_core.u_fifo_tx._0312_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0323_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0329_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0331_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0368_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1443_  (.A(\u_usb_host.u_core.u_fifo_tx._0316_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0342_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0345_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0350_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0369_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1444_  (.A(\u_usb_host.u_core.u_fifo_tx._0366_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0367_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0368_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0369_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0370_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1445_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0371_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1446_  (.A(\u_usb_host.u_core.u_fifo_tx._0317_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0326_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0346_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0348_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0372_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1447_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0371_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0372_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0373_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1448_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0374_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1449_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][6] ),
    .A2(net237),
    .A3(net197),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][6] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0375_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_fifo_tx._1450_  (.A(\u_usb_host.u_core.u_fifo_tx._0353_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0374_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0375_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0376_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1451_  (.A(\u_usb_host.u_core.u_fifo_tx._0365_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0370_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0373_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0376_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0377_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1452_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][6] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0360_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0377_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[6] ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1453_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[34][7] ),
    .B(net230),
    .C(net222),
    .X(\u_usb_host.u_core.u_fifo_tx._0378_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1454_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[58][7] ),
    .B(net257),
    .C(\u_usb_host.u_core.u_fifo_tx._0527_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0379_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1455_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[43][7] ),
    .B(net217),
    .C(net208),
    .X(\u_usb_host.u_core.u_fifo_tx._0380_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1456_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[8][7] ),
    .B(net239),
    .C(net211),
    .X(\u_usb_host.u_core.u_fifo_tx._0381_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1457_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[40][7] ),
    .B(net224),
    .C(net212),
    .X(\u_usb_host.u_core.u_fifo_tx._0382_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1458_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[50][7] ),
    .B(net250),
    .C(net229),
    .X(\u_usb_host.u_core.u_fifo_tx._0383_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1459_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[16][7] ),
    .B(net264),
    .C(net242),
    .X(\u_usb_host.u_core.u_fifo_tx._0384_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1460_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[57][7] ),
    .B(net254),
    .C(net233),
    .X(\u_usb_host.u_core.u_fifo_tx._0385_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1461_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[48][7] ),
    .B(net245),
    .C(net241),
    .X(\u_usb_host.u_core.u_fifo_tx._0386_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1462_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[18][7] ),
    .B(net262),
    .C(net231),
    .X(\u_usb_host.u_core.u_fifo_tx._0387_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1463_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[17][7] ),
    .B(net262),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0388_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1464_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[35][7] ),
    .B(net223),
    .C(net204),
    .X(\u_usb_host.u_core.u_fifo_tx._0389_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1465_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[59][7] ),
    .B(net249),
    .C(net209),
    .X(\u_usb_host.u_core.u_fifo_tx._0390_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1466_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[46][7] ),
    .B(net214),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0391_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1467_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[51][7] ),
    .B(net249),
    .C(net203),
    .X(\u_usb_host.u_core.u_fifo_tx._0392_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1468_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[49][7] ),
    .B(net244),
    .C(net205),
    .X(\u_usb_host.u_core.u_fifo_tx._0393_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1469_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[41][7] ),
    .B(net232),
    .C(net216),
    .X(\u_usb_host.u_core.u_fifo_tx._0394_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1470_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[33][7] ),
    .B(net220),
    .C(net207),
    .X(\u_usb_host.u_core.u_fifo_tx._0395_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1471_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[32][7] ),
    .B(net243),
    .C(net219),
    .X(\u_usb_host.u_core.u_fifo_tx._0396_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1472_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[63][7] ),
    .B(net272),
    .C(net254),
    .X(\u_usb_host.u_core.u_fifo_tx._0397_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1473_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[36][7] ),
    .B(net222),
    .C(net202),
    .X(\u_usb_host.u_core.u_fifo_tx._0398_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1474_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[37][7] ),
    .B(net224),
    .C(net191),
    .X(\u_usb_host.u_core.u_fifo_tx._0399_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1475_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[20][7] ),
    .B(net267),
    .C(net201),
    .X(\u_usb_host.u_core.u_fifo_tx._0400_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1476_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[14][7] ),
    .B(net234),
    .C(net186),
    .X(\u_usb_host.u_core.u_fifo_tx._0401_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1477_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[15][7] ),
    .B(net270),
    .C(net236),
    .X(\u_usb_host.u_core.u_fifo_tx._0402_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1478_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[28][7] ),
    .B(net259),
    .C(net196),
    .X(\u_usb_host.u_core.u_fifo_tx._0403_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1479_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[60][7] ),
    .B(net249),
    .C(net199),
    .X(\u_usb_host.u_core.u_fifo_tx._0404_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1480_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[47][7] ),
    .B(net269),
    .C(net214),
    .X(\u_usb_host.u_core.u_fifo_tx._0405_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1481_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[31][7] ),
    .B(net271),
    .C(net265),
    .X(\u_usb_host.u_core.u_fifo_tx._0406_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1482_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[61][7] ),
    .B(net250),
    .C(net195),
    .X(\u_usb_host.u_core.u_fifo_tx._0407_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1483_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[45][7] ),
    .B(net213),
    .C(net193),
    .X(\u_usb_host.u_core.u_fifo_tx._0408_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1484_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[38][7] ),
    .B(net224),
    .C(\u_usb_host.u_core.u_fifo_tx._0575_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0409_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1485_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[62][7] ),
    .B(net253),
    .C(net188),
    .X(\u_usb_host.u_core.u_fifo_tx._0410_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1486_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[52][7] ),
    .B(net246),
    .C(net200),
    .X(\u_usb_host.u_core.u_fifo_tx._0411_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1487_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[39][7] ),
    .B(\u_usb_host.u_core.u_fifo_tx._0504_ ),
    .C(net224),
    .X(\u_usb_host.u_core.u_fifo_tx._0412_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1488_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[53][7] ),
    .B(net250),
    .C(net190),
    .X(\u_usb_host.u_core.u_fifo_tx._0413_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1489_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[44][7] ),
    .B(net216),
    .C(net198),
    .X(\u_usb_host.u_core.u_fifo_tx._0414_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_fifo_tx._1490_  (.A(\u_usb_host.u_core.u_fifo_tx.ram[21][7] ),
    .B(net265),
    .C(net189),
    .X(\u_usb_host.u_core.u_fifo_tx._0415_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1491_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[19][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0546_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0559_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[26][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0416_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1492_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[13][7] ),
    .A2(net235),
    .A3(net194),
    .B1(\u_usb_host.u_core.u_fifo_tx._0393_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0401_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0417_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1493_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[5][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0572_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0576_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[6][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0418_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1494_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[3][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0545_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0553_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[1][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0419_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1495_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[27][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0533_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0577_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[4][7] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0418_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0420_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1496_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[2][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0543_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0578_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[7][7] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0419_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0421_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_fifo_tx._1497_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[25][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0521_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0526_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[24][7] ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0416_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0422_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_fifo_tx._1498_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[29][7] ),
    .A2(net260),
    .A3(net192),
    .B1(\u_usb_host.u_core.u_fifo_tx._0403_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0423_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_fifo_tx._1499_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[30][7] ),
    .A2(net261),
    .A3(net187),
    .B1(\u_usb_host.u_core.u_fifo_tx._0396_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0423_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0424_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1500_  (.A(\u_usb_host.u_core.u_fifo_tx._0420_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0421_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0422_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0424_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0425_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1501_  (.A(\u_usb_host.u_core.u_fifo_tx._0386_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0391_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0405_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0408_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0426_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1502_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[42][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0560_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0380_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0394_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0414_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0427_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1503_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[23][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0561_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0384_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0387_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0388_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0428_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1504_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[22][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0591_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0400_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0406_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0415_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0429_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1505_  (.A(\u_usb_host.u_core.u_fifo_tx._0426_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0427_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0428_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0429_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0430_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1506_  (.A(\u_usb_host.u_core.u_fifo_tx._0381_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0385_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0397_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0410_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0431_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1507_  (.A(\u_usb_host.u_core.u_fifo_tx._0379_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0390_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0404_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0407_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0432_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1508_  (.A(\u_usb_host.u_core.u_fifo_tx._0378_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0389_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0395_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0398_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0433_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1509_  (.A(\u_usb_host.u_core.u_fifo_tx._0382_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0399_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0409_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0412_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0434_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1510_  (.A(\u_usb_host.u_core.u_fifo_tx._0431_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0432_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0433_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0434_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0435_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1511_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[55][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0568_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0585_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[54][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0436_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1512_  (.A(\u_usb_host.u_core.u_fifo_tx._0383_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0392_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0411_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0413_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0437_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_fifo_tx._1513_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[56][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0537_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0436_ ),
    .C1(\u_usb_host.u_core.u_fifo_tx._0437_ ),
    .D1(\u_usb_host.u_core.u_fifo_tx._0518_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0438_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_fifo_tx._1514_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[10][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0528_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0538_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[9][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0439_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_fifo_tx._1515_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[12][7] ),
    .A2(net238),
    .A3(net196),
    .B1(\u_usb_host.u_core.u_fifo_tx._0536_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx.ram[11][7] ),
    .X(\u_usb_host.u_core.u_fifo_tx._0440_ ));
 sky130_fd_sc_hd__or4_2 \u_usb_host.u_core.u_fifo_tx._1516_  (.A(\u_usb_host.u_core.u_fifo_tx._0402_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0417_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0439_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0440_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0441_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_fifo_tx._1517_  (.A(\u_usb_host.u_core.u_fifo_tx._0430_ ),
    .B(\u_usb_host.u_core.u_fifo_tx._0435_ ),
    .C(\u_usb_host.u_core.u_fifo_tx._0438_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0441_ ),
    .X(\u_usb_host.u_core.u_fifo_tx._0442_ ));
 sky130_fd_sc_hd__o22a_2 \u_usb_host.u_core.u_fifo_tx._1518_  (.A1(\u_usb_host.u_core.u_fifo_tx.ram[0][7] ),
    .A2(\u_usb_host.u_core.u_fifo_tx._0519_ ),
    .B1(\u_usb_host.u_core.u_fifo_tx._0425_ ),
    .B2(\u_usb_host.u_core.u_fifo_tx._0442_ ),
    .X(\u_usb_host.u_core.fifo_tx_data_w[7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1519_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1520_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1521_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1522_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1523_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1524_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1525_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1526_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0752_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[24][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1527_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1528_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1529_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1530_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1531_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net488),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1532_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net479),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1533_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1534_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0783_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[55][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1535_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1536_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1537_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net501),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1538_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net492),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1539_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1540_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1541_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1542_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0751_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[23][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1543_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1544_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1545_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1546_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1547_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1548_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1549_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1550_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0750_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[22][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1551_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1552_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1553_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1554_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1555_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net488),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1556_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net479),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1557_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1558_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0782_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[54][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1559_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1560_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1561_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1562_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1563_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1564_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1565_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1566_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0749_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[21][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1567_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1568_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1569_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1570_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1571_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1572_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1573_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1574_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0781_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[53][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1575_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1576_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net513),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1577_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1578_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1579_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1580_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1581_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1582_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0748_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[20][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1583_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1584_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1585_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1586_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1587_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1588_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1589_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1590_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0747_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[19][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1591_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1592_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net513),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1593_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1594_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1595_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1596_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1597_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1598_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0780_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[52][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1599_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1600_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1601_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net501),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1602_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net492),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1603_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1604_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1605_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1606_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0746_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[18][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1607_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1608_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net516),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1609_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1610_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1611_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net488),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1612_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net479),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1613_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1614_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0779_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[51][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1615_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1616_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1617_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net501),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1618_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net492),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1619_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1620_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1621_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1622_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0745_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[17][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1623_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1624_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1625_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net501),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1626_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net492),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1627_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1628_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1629_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1630_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0744_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[16][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1631_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1632_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1633_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1634_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1635_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1636_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net479),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1637_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1638_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0778_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[50][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1639_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1640_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1641_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1642_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1643_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1644_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1645_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1646_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0743_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[15][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1647_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1648_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1649_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1650_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1651_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1652_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1653_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1654_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0777_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[49][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1655_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1656_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1657_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1658_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1659_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1660_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1661_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1662_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0742_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[14][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1663_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1664_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1665_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1666_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1667_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1668_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1669_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1670_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0741_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[13][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1671_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1672_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1673_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1674_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1675_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1676_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1677_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1678_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0776_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[48][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1679_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1680_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1681_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1682_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1683_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1684_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1685_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1686_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0740_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[12][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1687_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1688_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1689_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1690_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1691_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1692_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1693_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1694_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0775_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[47][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1695_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1696_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1697_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1698_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1699_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1700_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1701_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1702_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0739_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[11][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1703_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1704_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1705_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1706_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1707_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1708_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1709_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1710_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0738_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[10][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1711_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1712_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1713_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1714_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1715_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1716_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1717_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1718_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0774_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[46][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1719_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1720_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1721_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1722_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1723_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1724_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1725_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1726_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0737_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[9][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1727_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1728_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net509),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1729_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net501),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1730_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net492),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1731_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1732_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1733_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1734_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0773_ ),
    .D(net458),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[45][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1735_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1736_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1737_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net507),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1738_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1739_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1740_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1741_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1742_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0736_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[8][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1743_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1744_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1745_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1746_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1747_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1748_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1749_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1750_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0735_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[7][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1751_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1752_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1753_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1754_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1755_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1756_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1757_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1758_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0772_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[44][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1759_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1760_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1761_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1762_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1763_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1764_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1765_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1766_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0734_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[6][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1767_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1768_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1769_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1770_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1771_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1772_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1773_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1774_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0771_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[43][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1775_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1776_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1777_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1778_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1779_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1780_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1781_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1782_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0733_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[5][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1783_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1784_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1785_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1786_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1787_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1788_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1789_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1790_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0732_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[4][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1791_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1792_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1793_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1794_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1795_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1796_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1797_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1798_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0770_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[42][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1799_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1800_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1801_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1802_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1803_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1804_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1805_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1806_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0731_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[3][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1807_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1808_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1809_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1810_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1811_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1812_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1813_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1814_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0730_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[2][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1815_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net520),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1816_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1817_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1818_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1819_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1820_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net477),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1821_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1822_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0769_ ),
    .D(net460),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[41][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1823_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1824_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1825_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1826_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1827_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1828_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1829_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1830_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0729_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1831_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1832_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1833_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net507),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1834_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net498),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1835_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1836_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1837_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1838_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0768_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[40][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1839_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1840_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net513),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1841_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1842_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1843_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1844_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1845_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net469),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1846_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0728_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1847_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1848_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1849_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1850_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net498),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1851_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1852_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1853_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1854_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0767_ ),
    .D(net464),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[39][7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_tx._1855_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0000_ ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_tx._1856_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0001_ ),
    .RESET_B(net366),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1857_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0002_ ),
    .RESET_B(net367),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1858_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0003_ ),
    .RESET_B(net369),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1859_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0004_ ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1860_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0005_ ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1861_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0727_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0006_ ),
    .RESET_B(net377),
    .Q(\u_usb_host.u_core.u_fifo_tx.count[6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1862_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1863_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1864_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1865_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1866_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net490),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1867_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1868_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1869_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0766_ ),
    .D(net464),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[38][7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1870_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0007_ ),
    .RESET_B(net374),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1871_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0008_ ),
    .RESET_B(net374),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1872_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0009_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1873_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0010_ ),
    .RESET_B(net374),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1874_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0011_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._1875_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0726_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0012_ ),
    .RESET_B(net374),
    .Q(\u_usb_host.u_core.u_fifo_tx.rd_ptr[5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1876_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1877_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net516),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1878_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1879_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1880_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net490),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1881_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1882_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1883_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0765_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[37][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1884_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1885_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1886_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net507),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1887_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1888_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1889_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1890_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1891_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0721_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[63][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1892_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1893_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1894_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1895_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1896_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1897_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1898_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1899_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0764_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[36][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1900_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1901_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1902_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1903_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1904_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1905_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net481),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1906_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net473),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1907_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0763_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[35][7] ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1908_  (.CLK(clknet_leaf_3_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0019_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0721_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1909_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0020_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0722_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1910_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0021_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0723_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1911_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0022_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0724_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1912_  (.CLK(clknet_leaf_51_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0023_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0725_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1913_  (.CLK(clknet_leaf_3_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0024_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0726_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1914_  (.CLK(clknet_leaf_3_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0025_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0727_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1915_  (.CLK(clknet_leaf_54_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0026_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0728_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1916_  (.CLK(clknet_leaf_2_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0027_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0729_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1917_  (.CLK(clknet_leaf_51_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0028_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0730_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1918_  (.CLK(clknet_leaf_2_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0029_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0731_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1919_  (.CLK(clknet_leaf_53_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0030_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0732_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1920_  (.CLK(clknet_leaf_58_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0031_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0733_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1921_  (.CLK(clknet_leaf_58_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0032_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0734_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1922_  (.CLK(clknet_leaf_51_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0033_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0735_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1923_  (.CLK(clknet_leaf_4_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0034_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0736_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1924_  (.CLK(clknet_leaf_53_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0035_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0737_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1925_  (.CLK(clknet_leaf_53_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0036_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0738_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1926_  (.CLK(clknet_leaf_54_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0037_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0739_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1927_  (.CLK(clknet_leaf_55_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0038_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0740_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1928_  (.CLK(clknet_leaf_56_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0039_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0741_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1929_  (.CLK(clknet_leaf_55_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0040_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0742_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1930_  (.CLK(clknet_leaf_55_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0041_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0743_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1931_  (.CLK(clknet_leaf_44_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0042_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0744_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1932_  (.CLK(clknet_leaf_42_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0043_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0745_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1933_  (.CLK(clknet_leaf_42_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0044_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0746_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1934_  (.CLK(clknet_leaf_2_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0045_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0747_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1935_  (.CLK(clknet_leaf_54_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0046_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0748_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1936_  (.CLK(clknet_leaf_54_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0047_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0749_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1937_  (.CLK(clknet_leaf_44_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0048_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0750_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1938_  (.CLK(clknet_leaf_42_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0049_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0751_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1939_  (.CLK(clknet_leaf_51_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0050_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0752_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1940_  (.CLK(clknet_leaf_51_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0051_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0753_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1941_  (.CLK(clknet_3_0_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0052_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0754_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1942_  (.CLK(clknet_leaf_53_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0053_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0755_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1943_  (.CLK(clknet_leaf_56_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0054_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0756_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1944_  (.CLK(clknet_leaf_57_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0055_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0757_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1945_  (.CLK(clknet_leaf_57_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0056_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0758_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1946_  (.CLK(clknet_leaf_44_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0057_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0759_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1947_  (.CLK(clknet_leaf_53_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0058_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0760_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1948_  (.CLK(clknet_leaf_46_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0059_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0761_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1949_  (.CLK(clknet_leaf_38_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0060_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0762_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1950_  (.CLK(clknet_leaf_37_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0061_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0763_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1951_  (.CLK(clknet_leaf_38_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0062_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0764_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1952_  (.CLK(clknet_leaf_37_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0063_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0765_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1953_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0064_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0766_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1954_  (.CLK(clknet_leaf_37_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0065_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0767_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1955_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0066_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0768_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1956_  (.CLK(clknet_leaf_45_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0067_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0769_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1957_  (.CLK(clknet_leaf_45_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0068_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0770_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1958_  (.CLK(clknet_leaf_45_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0069_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0771_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1959_  (.CLK(clknet_leaf_45_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0070_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0772_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1960_  (.CLK(clknet_leaf_55_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0071_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0773_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1961_  (.CLK(clknet_leaf_43_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0072_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0774_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1962_  (.CLK(clknet_leaf_43_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0073_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0775_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1963_  (.CLK(clknet_leaf_43_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0074_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0776_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1964_  (.CLK(clknet_leaf_55_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0075_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0777_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1965_  (.CLK(clknet_leaf_46_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0076_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0778_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1966_  (.CLK(clknet_leaf_46_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0077_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0779_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1967_  (.CLK(clknet_leaf_46_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0078_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0780_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1968_  (.CLK(clknet_leaf_46_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0079_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0781_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1969_  (.CLK(clknet_3_3_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0080_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0782_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1970_  (.CLK(clknet_leaf_47_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0081_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0783_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1971_  (.CLK(clknet_leaf_47_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0082_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0784_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1972_  (.CLK(clknet_leaf_4_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0083_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0785_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1973_  (.CLK(clknet_leaf_49_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0084_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0786_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_fifo_tx._1974_  (.CLK(clknet_3_3_0_usb_clk),
    .GATE(\u_usb_host.u_core.u_fifo_tx._0085_ ),
    .GCLK(\u_usb_host.u_core.u_fifo_tx._0787_ ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1975_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1976_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net516),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1977_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1978_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1979_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1980_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1981_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1982_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0786_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[58][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1983_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1984_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net516),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1985_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1986_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1987_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net488),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1988_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1989_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1990_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0787_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[59][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1991_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1992_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1993_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1994_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1995_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1996_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net479),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1997_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1998_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0784_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[56][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._1999_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net523),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2000_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2001_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2002_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2003_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2004_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2005_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2006_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0785_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[57][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2007_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2008_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2009_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2010_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2011_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2012_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2013_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2014_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0758_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[30][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2015_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2016_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2017_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2018_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2019_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2020_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2021_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2022_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0760_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[32][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2023_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2024_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2025_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2026_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2027_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net486),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2028_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2029_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2030_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0754_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[26][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2031_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2032_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2033_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net502),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2034_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net493),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2035_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2036_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2037_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2038_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0755_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[27][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2039_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2040_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2041_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2042_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2043_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2044_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2045_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2046_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0756_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[28][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2047_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net517),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2048_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net510),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2049_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net500),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2050_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net491),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2051_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net484),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2052_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net474),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2053_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net466),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2054_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0757_ ),
    .D(net457),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[29][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2055_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net519),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2056_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net511),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2057_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net503),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2058_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net494),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2059_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net483),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2060_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net475),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2061_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net467),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2062_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0759_ ),
    .D(net459),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[31][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2063_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net518),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2064_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net512),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2065_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2066_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2067_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net485),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2068_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net476),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2069_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net468),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2070_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0753_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[25][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2071_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2072_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2073_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2074_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2075_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2076_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net481),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2077_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2078_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0762_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[34][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2079_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2080_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2081_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net505),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2082_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2083_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2084_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2085_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net471),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2086_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0761_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[33][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2087_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net521),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2088_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net516),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2089_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net504),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2090_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net495),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2091_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net487),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2092_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net478),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2093_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2094_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0724_ ),
    .D(net461),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[60][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2095_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net522),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2096_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net514),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2097_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net506),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2098_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net496),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2099_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net488),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2100_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net481),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2101_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net470),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2102_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0722_ ),
    .D(net462),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[61][7] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2103_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(\u_usb_host.u_core.u_fifo_tx.data_i[0] ),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][0] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2104_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net515),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][1] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2105_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net507),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][2] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2106_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net497),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][3] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2107_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net489),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][4] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2108_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net480),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][5] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2109_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net472),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][6] ));
 sky130_fd_sc_hd__dfxtp_1 \u_usb_host.u_core.u_fifo_tx._2110_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0723_ ),
    .D(net463),
    .Q(\u_usb_host.u_core.u_fifo_tx.ram[62][7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._2111_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0013_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._2112_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0014_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._2113_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0015_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._2114_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0016_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[3] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_fifo_tx._2115_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0017_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_fifo_tx._2116_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_fifo_tx._0725_ ),
    .D(\u_usb_host.u_core.u_fifo_tx._0018_ ),
    .RESET_B(net373),
    .Q(\u_usb_host.u_core.u_fifo_tx.wr_ptr[5] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._318_  (.A(net541),
    .Y(\u_usb_host.u_core.u_sie._081_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._319_  (.A(net543),
    .Y(\u_usb_host.u_core.u_sie._082_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._320_  (.A(net687),
    .Y(\u_usb_host.u_core.u_sie._083_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._321_  (.A(net540),
    .Y(\u_usb_host.u_core.u_sie._084_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._322_  (.A(\u_usb_host.u_core.status_rx_count_w[0] ),
    .Y(\u_usb_host.u_core.u_sie._085_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._323_  (.A(\u_usb_host.u_core.u_sie.in_transfer_q ),
    .Y(\u_usb_host.u_core.u_sie._086_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._324_  (.A(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .Y(\u_usb_host.u_core.u_sie._080_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._325_  (.A(\u_usb_host.u_core.u_sie.state_q[3] ),
    .B(\u_usb_host.u_core.u_sie.state_q[2] ),
    .Y(\u_usb_host.u_core.u_sie._087_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._326_  (.A(net542),
    .B(net543),
    .Y(\u_usb_host.u_core.u_sie._088_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._327_  (.A(\u_usb_host.u_core.u_sie._088_ ),
    .Y(\u_usb_host.u_core.u_sie._089_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_sie._328_  (.A(\u_usb_host.u_core.u_sie._087_ ),
    .B(\u_usb_host.u_core.u_sie._088_ ),
    .Y(\u_usb_host.u_core.u_sie._053_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._329_  (.A(\u_usb_host.u_core.u_sie._053_ ),
    .Y(\u_usb_host.u_core.status_sie_idle_w ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_sie._330_  (.A_N(\u_usb_host.u_core.u_sie.state_q[3] ),
    .B(\u_usb_host.u_core.u_sie.state_q[2] ),
    .Y(\u_usb_host.u_core.u_sie._090_ ));
 sky130_fd_sc_hd__or3_4 \u_usb_host.u_core.u_sie._331_  (.A(net541),
    .B(net425),
    .C(\u_usb_host.u_core.u_sie._090_ ),
    .X(\u_usb_host.u_core.u_sie._091_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._332_  (.A(\u_usb_host.u_core.u_sie._091_ ),
    .Y(\u_usb_host.u_core.u_sie._292_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._333_  (.A(\u_usb_host.u_core.u_sie.state_q[3] ),
    .B(\u_usb_host.u_core.u_sie.state_q[2] ),
    .Y(\u_usb_host.u_core.u_sie._092_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_sie._334_  (.A(\u_usb_host.u_core.u_sie.tx_ifs_q[1] ),
    .B(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ),
    .C(\u_usb_host.u_core.u_sie.tx_ifs_q[2] ),
    .X(\u_usb_host.u_core.u_sie._093_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._335_  (.A(\u_usb_host.u_core.u_sie.tx_ifs_q[3] ),
    .B(\u_usb_host.u_core.u_sie._093_ ),
    .X(\u_usb_host.u_core.u_sie._094_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._336_  (.A(\u_usb_host.u_core.u_sie.wait_eop_q ),
    .B(\u_usb_host.u_core.u_sie._094_ ),
    .Y(\u_usb_host.u_core.u_sie._095_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._337_  (.A(\u_usb_host.u_core.u_sie._095_ ),
    .Y(\u_usb_host.u_core.u_sie._096_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_sie._338_  (.A(net541),
    .B(\u_usb_host.u_core.u_sie._087_ ),
    .X(\u_usb_host.u_core.u_sie._097_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._339_  (.A(\u_usb_host.u_core.status_rx_count_w[13] ),
    .B(\u_usb_host.u_core.status_rx_count_w[12] ),
    .Y(\u_usb_host.u_core.u_sie._098_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._340_  (.A(\u_usb_host.u_core.status_rx_count_w[9] ),
    .B(\u_usb_host.u_core.status_rx_count_w[8] ),
    .Y(\u_usb_host.u_core.u_sie._099_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._341_  (.A(\u_usb_host.u_core.status_rx_count_w[9] ),
    .B(\u_usb_host.u_core.status_rx_count_w[8] ),
    .C(\u_usb_host.u_core.status_rx_count_w[11] ),
    .D(\u_usb_host.u_core.status_rx_count_w[10] ),
    .X(\u_usb_host.u_core.u_sie._100_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._342_  (.A(\u_usb_host.u_core.status_rx_count_w[5] ),
    .B(\u_usb_host.u_core.status_rx_count_w[4] ),
    .Y(\u_usb_host.u_core.u_sie._101_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._343_  (.A(\u_usb_host.u_core.status_rx_count_w[5] ),
    .B(\u_usb_host.u_core.status_rx_count_w[4] ),
    .C(\u_usb_host.u_core.status_rx_count_w[7] ),
    .D(\u_usb_host.u_core.status_rx_count_w[6] ),
    .X(\u_usb_host.u_core.u_sie._102_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_sie._344_  (.A(\u_usb_host.u_core.transfer_start_q ),
    .B(net114),
    .Y(\u_usb_host.u_core.u_sie._103_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._345_  (.A(\u_usb_host.u_core.u_sie._103_ ),
    .Y(\u_usb_host.u_core.u_sie._070_ ));
 sky130_fd_sc_hd__nand2b_2 \u_usb_host.u_core.u_sie._346_  (.A_N(\u_usb_host.u_core.u_sie.state_q[2] ),
    .B(\u_usb_host.u_core.u_sie.state_q[3] ),
    .Y(\u_usb_host.u_core.u_sie._104_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._347_  (.A(net541),
    .B(\u_usb_host.u_core.u_sie._104_ ),
    .Y(\u_usb_host.u_core.u_sie._105_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._348_  (.A(net541),
    .B(\u_usb_host.u_core.u_sie._104_ ),
    .X(\u_usb_host.u_core.u_sie._106_ ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._349_  (.A(net543),
    .B(\u_usb_host.u_core.u_sie._106_ ),
    .Y(\u_usb_host.u_core.u_sie._107_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._350_  (.A(net425),
    .B(\u_usb_host.u_core.u_sie._105_ ),
    .Y(\u_usb_host.u_core.u_sie._108_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core.u_sie._351_  (.A1(\u_usb_host.u_core.u_sie._086_ ),
    .A2(\u_usb_host.u_core.u_sie.send_sof_q ),
    .B1(\u_usb_host.u_core.u_sie._107_ ),
    .C1(net540),
    .X(\u_usb_host.u_core.u_sie._109_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._352_  (.A(net543),
    .B(\u_usb_host.u_core.u_sie._090_ ),
    .Y(\u_usb_host.u_core.u_sie._110_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._353_  (.A1(net543),
    .A2(\u_usb_host.u_core.u_sie.utmi_txready_i ),
    .B1(\u_usb_host.u_core.u_sie._090_ ),
    .X(\u_usb_host.u_core.u_sie._111_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._354_  (.A(\u_usb_host.u_core.status_rx_count_w[0] ),
    .B(\u_usb_host.u_core.status_rx_count_w[3] ),
    .C(\u_usb_host.u_core.status_rx_count_w[2] ),
    .D(\u_usb_host.u_core.status_rx_count_w[15] ),
    .X(\u_usb_host.u_core.u_sie._112_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._355_  (.A(\u_usb_host.u_core.status_rx_count_w[1] ),
    .B(\u_usb_host.u_core.status_rx_count_w[13] ),
    .C(\u_usb_host.u_core.status_rx_count_w[12] ),
    .D(\u_usb_host.u_core.status_rx_count_w[14] ),
    .X(\u_usb_host.u_core.u_sie._113_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_core.u_sie._356_  (.A(\u_usb_host.u_core.u_sie._089_ ),
    .B(\u_usb_host.u_core.u_sie._092_ ),
    .C(\u_usb_host.u_core.u_sie._095_ ),
    .Y(\u_usb_host.u_core.u_sie._114_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._357_  (.A(net425),
    .B(\u_usb_host.u_core.u_sie._092_ ),
    .Y(\u_usb_host.u_core.u_sie._115_ ));
 sky130_fd_sc_hd__nand2_2 \u_usb_host.u_core.u_sie._358_  (.A(\u_usb_host.u_core.u_sie._081_ ),
    .B(\u_usb_host.u_core.u_sie._110_ ),
    .Y(\u_usb_host.u_core.u_sie._116_ ));
 sky130_fd_sc_hd__and2_2 \u_usb_host.u_core.u_sie._359_  (.A(net541),
    .B(\u_usb_host.u_core.u_sie._110_ ),
    .X(\u_usb_host.u_core.u_sie._117_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_core.u_sie._360_  (.A1(\u_usb_host.u_core.u_sie._088_ ),
    .A2(\u_usb_host.u_core.u_sie._092_ ),
    .B1(\u_usb_host.u_core.u_sie._103_ ),
    .C1(\u_usb_host.u_core.u_sie._111_ ),
    .X(\u_usb_host.u_core.u_sie._118_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._361_  (.A(\u_usb_host.u_core.u_sie._100_ ),
    .B(\u_usb_host.u_core.u_sie._102_ ),
    .C(\u_usb_host.u_core.u_sie._112_ ),
    .D(\u_usb_host.u_core.u_sie._113_ ),
    .X(\u_usb_host.u_core.u_sie._119_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_sie._362_  (.A_N(\u_usb_host.u_core.u_sie.state_q[3] ),
    .B_N(\u_usb_host.u_core.u_sie.state_q[2] ),
    .C(net542),
    .D(\u_usb_host.u_core.u_sie.utmi_txready_i ),
    .X(\u_usb_host.u_core.u_sie._120_ ));
 sky130_fd_sc_hd__nand2_4 \u_usb_host.u_core.u_sie._363_  (.A(net540),
    .B(\u_usb_host.u_core.u_sie._097_ ),
    .Y(\u_usb_host.u_core.u_sie._121_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._364_  (.A(\u_usb_host.u_core.u_sie._119_ ),
    .B(\u_usb_host.u_core.u_sie._121_ ),
    .Y(\u_usb_host.u_core.u_sie._122_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core.u_sie._365_  (.A(\u_usb_host.u_core.u_sie._109_ ),
    .B(\u_usb_host.u_core.u_sie._114_ ),
    .C(\u_usb_host.u_core.u_sie._122_ ),
    .D_N(\u_usb_host.u_core.u_sie._118_ ),
    .X(\u_usb_host.u_core.u_sie.next_state_r[2] ));
 sky130_fd_sc_hd__nor3_4 \u_usb_host.u_core.u_sie._366_  (.A(\u_usb_host.u_core.u_sie._081_ ),
    .B(net425),
    .C(\u_usb_host.u_core.u_sie._104_ ),
    .Y(\u_usb_host.u_core.u_sie._123_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._367_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[1] ),
    .B(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ),
    .C(\u_usb_host.u_core.u_sie.last_tx_time_q[2] ),
    .X(\u_usb_host.u_core.u_sie._124_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._368_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[3] ),
    .B(\u_usb_host.u_core.u_sie._124_ ),
    .X(\u_usb_host.u_core.u_sie._125_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._369_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[3] ),
    .B(\u_usb_host.u_core.u_sie.last_tx_time_q[4] ),
    .C(\u_usb_host.u_core.u_sie._124_ ),
    .X(\u_usb_host.u_core.u_sie._126_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._370_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[5] ),
    .B(\u_usb_host.u_core.u_sie.last_tx_time_q[4] ),
    .C(\u_usb_host.u_core.u_sie._125_ ),
    .X(\u_usb_host.u_core.u_sie._127_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._371_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[6] ),
    .B(\u_usb_host.u_core.u_sie._127_ ),
    .X(\u_usb_host.u_core.u_sie._128_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._372_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[7] ),
    .B(\u_usb_host.u_core.u_sie.last_tx_time_q[6] ),
    .C(\u_usb_host.u_core.u_sie._127_ ),
    .X(\u_usb_host.u_core.u_sie._129_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._373_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[8] ),
    .B(\u_usb_host.u_core.u_sie._129_ ),
    .X(\u_usb_host.u_core.u_sie._130_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._374_  (.A(\u_usb_host.u_core.u_sie.wait_resp_q ),
    .B(\u_usb_host.u_core.u_sie._130_ ),
    .Y(\u_usb_host.u_core.u_sie._131_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._375_  (.A1(\u_usb_host.u_core.u_sie._084_ ),
    .A2(\u_usb_host.u_core.u_sie._119_ ),
    .B1(\u_usb_host.u_core.u_sie._097_ ),
    .X(\u_usb_host.u_core.u_sie._132_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._376_  (.A(\u_usb_host.u_core.u_sie.data_ready_w ),
    .B(\u_usb_host.u_core.u_sie._123_ ),
    .Y(\u_usb_host.u_core.u_sie._133_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._377_  (.A(net543),
    .B(\u_usb_host.u_core.u_sie._084_ ),
    .C(\u_usb_host.u_core.u_sie._105_ ),
    .X(\u_usb_host.u_core.u_sie._134_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._378_  (.A1(\u_usb_host.u_core.u_sie.wait_resp_q ),
    .A2(\u_usb_host.u_core.u_sie._084_ ),
    .B1(\u_usb_host.u_core.u_sie._292_ ),
    .X(\u_usb_host.u_core.u_sie._135_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._379_  (.A(\u_usb_host.u_core.u_sie._081_ ),
    .B(net543),
    .C(\u_usb_host.u_core.u_sie._087_ ),
    .X(\u_usb_host.u_core.u_sie._136_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_core.u_sie._380_  (.A(net541),
    .B(net425),
    .C_N(\u_usb_host.u_core.u_sie._087_ ),
    .X(\u_usb_host.u_core.u_sie._137_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_sie._381_  (.A_N(\u_usb_host.u_core.u_sie.send_sof_q ),
    .B(\u_usb_host.u_core.u_sie._107_ ),
    .C(net540),
    .D(\u_usb_host.u_core.u_sie.in_transfer_q ),
    .X(\u_usb_host.u_core.u_sie._138_ ));
 sky130_fd_sc_hd__nor3_4 \u_usb_host.u_core.u_sie._382_  (.A(\u_usb_host.u_core.u_sie._081_ ),
    .B(net425),
    .C(\u_usb_host.u_core.u_sie._090_ ),
    .Y(\u_usb_host.u_core.u_sie._139_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._383_  (.A(\u_usb_host.u_core.u_sie.state_q[0] ),
    .B(\u_usb_host.u_core.u_sie._104_ ),
    .Y(\u_usb_host.u_core.u_sie._140_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._384_  (.A1(\u_usb_host.u_core.u_sie._084_ ),
    .A2(\u_usb_host.u_core.u_sie._139_ ),
    .B1(\u_usb_host.u_core.u_sie._138_ ),
    .C1(\u_usb_host.u_core.u_sie._132_ ),
    .X(\u_usb_host.u_core.u_sie._141_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._385_  (.A1(net543),
    .A2(net540),
    .B1(\u_usb_host.u_core.u_sie._141_ ),
    .X(\u_usb_host.u_core.u_sie._142_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_sie._386_  (.A1(net543),
    .A2(net540),
    .B1(\u_usb_host.u_core.u_sie._110_ ),
    .B2(\u_usb_host.u_core.u_sie._115_ ),
    .X(\u_usb_host.u_core.u_sie._143_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_sie._387_  (.A1(net541),
    .A2(\u_usb_host.u_core.u_sie._095_ ),
    .A3(\u_usb_host.u_core.u_sie._140_ ),
    .B1(\u_usb_host.u_core.u_sie._134_ ),
    .X(\u_usb_host.u_core.u_sie._144_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._388_  (.A1(\u_usb_host.u_core.u_sie.rx_active_q[0] ),
    .A2(\u_usb_host.u_core.u_sie._136_ ),
    .B1(\u_usb_host.u_core.u_sie._143_ ),
    .C1(\u_usb_host.u_core.u_sie._144_ ),
    .X(\u_usb_host.u_core.u_sie._145_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core.u_sie._389_  (.A(\u_usb_host.u_core.u_sie._135_ ),
    .B(\u_usb_host.u_core.u_sie._145_ ),
    .C(\u_usb_host.u_core.u_sie._142_ ),
    .D_N(\u_usb_host.u_core.u_sie._133_ ),
    .X(\u_usb_host.u_core.u_sie._146_ ));
 sky130_fd_sc_hd__and3_2 \u_usb_host.u_core.u_sie._390_  (.A(net541),
    .B(net543),
    .C(\u_usb_host.u_core.u_sie._087_ ),
    .X(\u_usb_host.u_core.u_sie._147_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._391_  (.A(\u_usb_host.u_core.u_sie._147_ ),
    .Y(\u_usb_host.u_core.u_sie._148_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._392_  (.A1(\u_usb_host.u_core.u_sie._123_ ),
    .A2(\u_usb_host.u_core.u_sie._131_ ),
    .B1(\u_usb_host.u_core.u_sie._146_ ),
    .X(\u_usb_host.u_core.u_sie.next_state_r[0] ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._393_  (.A(\u_usb_host.u_core.u_sie._083_ ),
    .B(\u_usb_host.u_core.u_sie._123_ ),
    .X(\u_usb_host.u_core.u_sie._149_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._394_  (.A(\u_usb_host.u_core.status_response_w[3] ),
    .B(\u_usb_host.u_core.status_response_w[7] ),
    .Y(\u_usb_host.u_core.u_sie._150_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._395_  (.A(\u_usb_host.u_core.status_response_w[3] ),
    .B(\u_usb_host.u_core.status_response_w[7] ),
    .Y(\u_usb_host.u_core.u_sie._151_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core.u_sie._396_  (.A(\u_usb_host.u_core.status_response_w[2] ),
    .B(\u_usb_host.u_core.status_response_w[5] ),
    .C(\u_usb_host.u_core.status_response_w[4] ),
    .D_N(\u_usb_host.u_core.status_response_w[6] ),
    .X(\u_usb_host.u_core.u_sie._152_ ));
 sky130_fd_sc_hd__and4bb_1 \u_usb_host.u_core.u_sie._397_  (.A_N(\u_usb_host.u_core.u_sie._150_ ),
    .B_N(\u_usb_host.u_core.u_sie._152_ ),
    .C(\u_usb_host.u_core.u_sie._151_ ),
    .D(\u_usb_host.u_core.status_response_w[0] ),
    .X(\u_usb_host.u_core.u_sie._153_ ));
 sky130_fd_sc_hd__and4b_1 \u_usb_host.u_core.u_sie._398_  (.A_N(\u_usb_host.u_core.u_sie.rx_active_q[0] ),
    .B(\u_usb_host.u_core.status_response_w[1] ),
    .C(\u_usb_host.u_core.u_sie._136_ ),
    .D(\u_usb_host.u_core.u_sie._153_ ),
    .X(\u_usb_host.u_core.u_sie._154_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._399_  (.A(\u_usb_host.u_core.u_sie.send_ack_q ),
    .B(\u_usb_host.u_core.u_sie._154_ ),
    .Y(\u_usb_host.u_core.u_sie._155_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._400_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[5] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[4] ),
    .C(\u_usb_host.u_core.u_sie.crc_sum_q[6] ),
    .D(\u_usb_host.u_core.u_sie.crc_sum_q[7] ),
    .X(\u_usb_host.u_core.u_sie._156_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core.u_sie._401_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[1] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .C(\u_usb_host.u_core.u_sie.crc_sum_q[2] ),
    .D_N(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .X(\u_usb_host.u_core.u_sie._157_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._402_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[12] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[15] ),
    .Y(\u_usb_host.u_core.u_sie._158_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._403_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[9] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[8] ),
    .C(\u_usb_host.u_core.u_sie.crc_sum_q[11] ),
    .D(\u_usb_host.u_core.u_sie.crc_sum_q[10] ),
    .X(\u_usb_host.u_core.u_sie._159_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_core.u_sie._404_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[14] ),
    .B(\u_usb_host.u_core.u_sie._158_ ),
    .C(\u_usb_host.u_core.u_sie._159_ ),
    .D_N(\u_usb_host.u_core.u_sie.crc_sum_q[13] ),
    .X(\u_usb_host.u_core.u_sie._160_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_core.u_sie._405_  (.A1(\u_usb_host.u_core.u_sie._156_ ),
    .A2(\u_usb_host.u_core.u_sie._157_ ),
    .A3(\u_usb_host.u_core.u_sie._160_ ),
    .B1(\u_usb_host.u_core.u_sie._154_ ),
    .C1(\u_usb_host.u_core.u_sie.in_transfer_q ),
    .X(\u_usb_host.u_core.u_sie._043_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_sie._406_  (.A1_N(\u_usb_host.u_core.u_sie._155_ ),
    .A2_N(\u_usb_host.u_core.u_sie._043_ ),
    .B1(net540),
    .B2(\u_usb_host.u_core.u_sie._135_ ),
    .X(\u_usb_host.u_core.u_sie._161_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_sie._407_  (.A1(net542),
    .A2(\u_usb_host.u_core.u_sie._131_ ),
    .A3(\u_usb_host.u_core.u_sie._149_ ),
    .B1(\u_usb_host.u_core.u_sie._161_ ),
    .X(\u_usb_host.u_core.u_sie._162_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_sie._408_  (.A1(\u_usb_host.u_core.u_sie.state_q[3] ),
    .A2(\u_usb_host.u_core.u_sie.state_q[2] ),
    .A3(\u_usb_host.u_core.u_sie._089_ ),
    .B1(\u_usb_host.u_core.u_sie._134_ ),
    .C1(\u_usb_host.u_core.u_sie._140_ ),
    .X(\u_usb_host.u_core.u_sie._163_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_core.u_sie._409_  (.A1(net540),
    .A2(\u_usb_host.u_core.u_sie._139_ ),
    .B1(\u_usb_host.u_core.u_sie._162_ ),
    .C1(\u_usb_host.u_core.u_sie._163_ ),
    .D1(\u_usb_host.u_core.u_sie._114_ ),
    .X(\u_usb_host.u_core.u_sie.next_state_r[3] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._410_  (.A(net525),
    .B(\u_usb_host.u_core.u_sie._103_ ),
    .Y(\u_usb_host.u_core.u_sie._164_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._411_  (.A(\u_usb_host.u_core.u_sie.data_ready_w ),
    .B(\u_usb_host.u_core.u_sie._137_ ),
    .Y(\u_usb_host.u_core.u_sie._165_ ));
 sky130_fd_sc_hd__o2bb2a_1 \u_usb_host.u_core.u_sie._412_  (.A1_N(\u_usb_host.u_core.u_sie.rx_active_q[0] ),
    .A2_N(\u_usb_host.u_core.u_sie._136_ ),
    .B1(net106),
    .B2(\u_usb_host.u_core.u_sie._165_ ),
    .X(\u_usb_host.u_core.u_sie._076_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_core.u_sie._413_  (.A(net541),
    .B(net540),
    .C(\u_usb_host.u_core.u_sie._110_ ),
    .X(\u_usb_host.u_core.u_sie._042_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._414_  (.A(net113),
    .B(\u_usb_host.u_core.u_sie._042_ ),
    .X(\u_usb_host.u_core.u_sie._077_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._415_  (.A(\u_usb_host.u_core.u_sie._103_ ),
    .B(\u_usb_host.u_core.u_sie._133_ ),
    .Y(\u_usb_host.u_core.u_sie._071_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._416_  (.A(\u_usb_host.u_core.u_sie._123_ ),
    .B(net106),
    .Y(\u_usb_host.u_core.u_sie._166_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_core.u_sie._417_  (.A1(\u_usb_host.u_core.u_sie._083_ ),
    .A2(\u_usb_host.u_core.u_sie.crc_byte_w ),
    .A3(\u_usb_host.u_core.u_sie._137_ ),
    .B1(net101),
    .C1(\u_usb_host.u_core.u_sie._121_ ),
    .X(\u_usb_host.u_core.u_sie._167_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._418_  (.A(\u_usb_host.u_core.u_sie._122_ ),
    .B(\u_usb_host.u_core.u_sie._167_ ),
    .Y(\u_usb_host.u_core.u_sie._069_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._419_  (.A1(\u_usb_host.u_core.u_sie.state_q[2] ),
    .A2(net542),
    .B1(\u_usb_host.u_core.u_sie.state_q[3] ),
    .X(\u_usb_host.u_core.u_sie._168_ ));
 sky130_fd_sc_hd__a21oi_4 \u_usb_host.u_core.u_sie._420_  (.A1(\u_usb_host.u_core.u_sie._081_ ),
    .A2(\u_usb_host.u_core.u_sie._087_ ),
    .B1(\u_usb_host.u_core.u_sie._168_ ),
    .Y(\u_usb_host.u_core.u_sie.utmi_txvalid_o ));
 sky130_fd_sc_hd__a21oi_4 \u_usb_host.u_core.u_sie._421_  (.A1(net584),
    .A2(\u_usb_host.u_core.u_sie.utmi_txvalid_o ),
    .B1(net114),
    .Y(\u_usb_host.u_core.u_sie._169_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._422_  (.A(\u_usb_host.u_core.u_sie._130_ ),
    .B(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._068_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._423_  (.A(\u_usb_host.u_core.u_sie._135_ ),
    .B(\u_usb_host.u_core.u_sie._136_ ),
    .Y(\u_usb_host.u_core.u_sie._072_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._424_  (.A1(\u_usb_host.u_core.u_sie._087_ ),
    .A2(\u_usb_host.u_core.u_sie._089_ ),
    .B1(\u_usb_host.u_core.u_sie._123_ ),
    .X(\u_usb_host.u_core.u_sie._170_ ));
 sky130_fd_sc_hd__o221a_1 \u_usb_host.u_core.u_sie._425_  (.A1(\u_usb_host.u_core.u_sie.data_ready_w ),
    .A2(net183),
    .B1(\u_usb_host.u_core.u_sie._148_ ),
    .B2(net540),
    .C1(\u_usb_host.u_core.u_sie._170_ ),
    .X(\u_usb_host.u_core.u_sie._078_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._426_  (.A1(net542),
    .A2(\u_usb_host.u_core.u_sie._131_ ),
    .B1(net101),
    .Y(\u_usb_host.u_core.u_sie._074_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._427_  (.A1(\u_usb_host.u_core.u_sie._123_ ),
    .A2(net106),
    .B1(\u_usb_host.u_core.u_sie._071_ ),
    .X(\u_usb_host.u_core.u_sie._075_ ));
 sky130_fd_sc_hd__o21ai_2 \u_usb_host.u_core.u_sie._428_  (.A1(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .A2(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .B1(net581),
    .Y(\u_usb_host.u_core.u_sie._063_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_core.u_sie._429_  (.A_N(\u_usb_host.u_core.u_sie.wait_eop_q ),
    .B(\u_usb_host.u_core.u_sie._063_ ),
    .Y(\u_usb_host.u_core.u_sie._171_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._430_  (.A(\u_usb_host.u_core.u_sie._094_ ),
    .B(\u_usb_host.u_core.u_sie._171_ ),
    .X(\u_usb_host.u_core.u_sie._067_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._431_  (.A(\u_usb_host.u_core.u_sie.send_sof_q ),
    .B(\u_usb_host.u_core.u_sie._092_ ),
    .Y(\u_usb_host.u_core.u_sie._172_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_sie._432_  (.A1(net542),
    .A2(\u_usb_host.u_core.u_sie._096_ ),
    .A3(\u_usb_host.u_core.u_sie._140_ ),
    .B1(\u_usb_host.u_core.u_sie._117_ ),
    .C1(\u_usb_host.u_core.u_sie._070_ ),
    .X(\u_usb_host.u_core.u_sie._173_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_sie._433_  (.A1(\u_usb_host.u_core.u_sie._088_ ),
    .A2(\u_usb_host.u_core.u_sie._095_ ),
    .A3(\u_usb_host.u_core.u_sie._172_ ),
    .B1(\u_usb_host.u_core.u_sie._173_ ),
    .C1(\u_usb_host.u_core.u_sie._141_ ),
    .X(\u_usb_host.u_core.u_sie._174_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_core.u_sie._434_  (.A1(\u_usb_host.u_core.u_sie.state_q[3] ),
    .A2(\u_usb_host.u_core.u_sie.state_q[2] ),
    .A3(net542),
    .B1(\u_usb_host.u_core.u_sie._162_ ),
    .C1(\u_usb_host.u_core.u_sie._174_ ),
    .X(\u_usb_host.u_core.u_sie.next_state_r[1] ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._435_  (.A1(\u_usb_host.u_core.u_sie._091_ ),
    .A2(\u_usb_host.u_core.u_sie._106_ ),
    .B1(\u_usb_host.u_core.u_sie._084_ ),
    .X(\u_usb_host.u_core.u_sie._175_ ));
 sky130_fd_sc_hd__o211ai_1 \u_usb_host.u_core.u_sie._436_  (.A1(\u_usb_host.u_core.u_sie._080_ ),
    .A2(\u_usb_host.u_core.u_sie.rx_active_q[3] ),
    .B1(\u_usb_host.u_core.u_sie._063_ ),
    .C1(\u_usb_host.u_core.u_sie._175_ ),
    .Y(\u_usb_host.u_core.u_sie._066_ ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_core.u_sie._437_  (.A(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .B(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .C(\u_usb_host.u_core.u_sie.utmi_linestate_q[1] ),
    .D(\u_usb_host.u_core.u_sie.utmi_linestate_q[0] ),
    .Y(\u_usb_host.u_core.u_sie.se0_detect_w ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._438_  (.A(\u_usb_host.u_core.resp_expected_q ),
    .B(\u_usb_host.u_core.in_transfer_q ),
    .X(\u_usb_host.u_core.u_sie._079_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._439_  (.A(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .B(net574),
    .X(\u_usb_host.u_core.u_sie._065_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._440_  (.A(\u_usb_host.u_core.u_sie._080_ ),
    .B(\u_usb_host.u_core.u_sie.utmi_rxvalid_i ),
    .X(\u_usb_host.u_core.u_sie.shift_en_w ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_core.u_sie._441_  (.A(\u_usb_host.u_core.u_sie._082_ ),
    .B(\u_usb_host.u_core.u_sie._121_ ),
    .Y(\u_usb_host.u_core.fifo_tx_pop_w ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._442_  (.A(\u_usb_host.u_core.u_sie.crc5_out_w[0] ),
    .B(net113),
    .Y(\u_usb_host.u_core.u_sie._054_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._443_  (.A(\u_usb_host.u_core.u_sie.crc5_out_w[1] ),
    .B(net113),
    .Y(\u_usb_host.u_core.u_sie._055_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._444_  (.A(\u_usb_host.u_core.u_sie.crc5_out_w[2] ),
    .B(net113),
    .Y(\u_usb_host.u_core.u_sie._056_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._445_  (.A(\u_usb_host.u_core.u_sie.crc5_out_w[3] ),
    .B(net113),
    .Y(\u_usb_host.u_core.u_sie._057_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._446_  (.A(\u_usb_host.u_core.u_sie.crc5_out_w[4] ),
    .B(net114),
    .Y(\u_usb_host.u_core.u_sie._058_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._447_  (.A1(net425),
    .A2(\u_usb_host.u_core.u_sie._097_ ),
    .B1(\u_usb_host.u_core.u_sie._123_ ),
    .X(\u_usb_host.u_core.u_sie._176_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._448_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[0] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._016_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._449_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[1] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._023_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._450_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[2] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._024_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._451_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[3] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._025_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._452_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[4] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._026_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._453_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[5] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._027_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._454_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[6] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._028_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._455_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[7] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._029_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._456_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[8] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._030_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._457_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[9] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._031_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._458_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[10] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._017_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._459_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[11] ),
    .B(net112),
    .X(\u_usb_host.u_core.u_sie._018_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._460_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[12] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._019_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._461_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[13] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._020_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._462_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[14] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._021_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._463_  (.A(\u_usb_host.u_core.u_sie.crc_out_w[15] ),
    .B(net111),
    .X(\u_usb_host.u_core.u_sie._022_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._464_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[0] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._044_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._465_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[1] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._045_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._466_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[2] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._046_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._467_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[3] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._047_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._468_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[4] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._048_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._469_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[5] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._049_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._470_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[6] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._050_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._471_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[7] ),
    .B(\u_usb_host.u_core.u_sie._053_ ),
    .X(\u_usb_host.u_core.u_sie._051_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._472_  (.A(\u_usb_host.u_core.resp_expected_q ),
    .B(\u_usb_host.u_core.u_sie._133_ ),
    .X(\u_usb_host.u_core.u_sie._064_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._473_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[0] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._085_ ),
    .X(\u_usb_host.u_core.u_sie._000_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._474_  (.A(\u_usb_host.u_core.status_rx_count_w[1] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._177_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._475_  (.A(\u_usb_host.u_core.status_rx_count_w[1] ),
    .B(net422),
    .X(\u_usb_host.u_core.u_sie._178_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_sie._476_  (.A(\u_usb_host.u_core.status_rx_count_w[0] ),
    .B(\u_usb_host.u_core.u_sie._177_ ),
    .C(\u_usb_host.u_core.u_sie._178_ ),
    .Y(\u_usb_host.u_core.u_sie._179_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._477_  (.A1(\u_usb_host.u_core.u_sie._177_ ),
    .A2(\u_usb_host.u_core.u_sie._178_ ),
    .B1(\u_usb_host.u_core.status_rx_count_w[0] ),
    .X(\u_usb_host.u_core.u_sie._180_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._478_  (.A1(net100),
    .A2(\u_usb_host.u_core.u_sie._179_ ),
    .A3(\u_usb_host.u_core.u_sie._180_ ),
    .B1(net105),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[1] ),
    .X(\u_usb_host.u_core.u_sie._007_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._479_  (.A(\u_usb_host.u_core.status_rx_count_w[2] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._181_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._480_  (.A(\u_usb_host.u_core.status_rx_count_w[2] ),
    .B(net422),
    .X(\u_usb_host.u_core.u_sie._182_ ));
 sky130_fd_sc_hd__a21boi_1 \u_usb_host.u_core.u_sie._481_  (.A1(\u_usb_host.u_core.status_rx_count_w[0] ),
    .A2(\u_usb_host.u_core.u_sie._178_ ),
    .B1_N(\u_usb_host.u_core.u_sie._177_ ),
    .Y(\u_usb_host.u_core.u_sie._183_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_sie._482_  (.A(\u_usb_host.u_core.u_sie._181_ ),
    .B(\u_usb_host.u_core.u_sie._182_ ),
    .C(\u_usb_host.u_core.u_sie._183_ ),
    .X(\u_usb_host.u_core.u_sie._184_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._483_  (.A1(\u_usb_host.u_core.u_sie._181_ ),
    .A2(\u_usb_host.u_core.u_sie._182_ ),
    .B1(\u_usb_host.u_core.u_sie._183_ ),
    .Y(\u_usb_host.u_core.u_sie._185_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._484_  (.A1(net100),
    .A2(\u_usb_host.u_core.u_sie._184_ ),
    .A3(\u_usb_host.u_core.u_sie._185_ ),
    .B1(net105),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[2] ),
    .X(\u_usb_host.u_core.u_sie._008_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_core.u_sie._485_  (.A_N(\u_usb_host.u_core.u_sie._182_ ),
    .B(\u_usb_host.u_core.u_sie._184_ ),
    .Y(\u_usb_host.u_core.u_sie._186_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._486_  (.A(\u_usb_host.u_core.status_rx_count_w[3] ),
    .B(net424),
    .Y(\u_usb_host.u_core.u_sie._187_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._487_  (.A(\u_usb_host.u_core.status_rx_count_w[3] ),
    .B(net424),
    .X(\u_usb_host.u_core.u_sie._188_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._488_  (.A(\u_usb_host.u_core.u_sie._187_ ),
    .B(\u_usb_host.u_core.u_sie._188_ ),
    .X(\u_usb_host.u_core.u_sie._189_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._489_  (.A(\u_usb_host.u_core.u_sie._186_ ),
    .B(\u_usb_host.u_core.u_sie._189_ ),
    .Y(\u_usb_host.u_core.u_sie._190_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._490_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[3] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._190_ ),
    .X(\u_usb_host.u_core.u_sie._009_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._491_  (.A1(\u_usb_host.u_core.status_rx_count_w[3] ),
    .A2(\u_usb_host.u_core.status_rx_count_w[2] ),
    .B1(net424),
    .Y(\u_usb_host.u_core.u_sie._191_ ));
 sky130_fd_sc_hd__o41a_1 \u_usb_host.u_core.u_sie._492_  (.A1(\u_usb_host.u_core.u_sie._181_ ),
    .A2(\u_usb_host.u_core.u_sie._182_ ),
    .A3(\u_usb_host.u_core.u_sie._183_ ),
    .A4(\u_usb_host.u_core.u_sie._187_ ),
    .B1(\u_usb_host.u_core.u_sie._191_ ),
    .X(\u_usb_host.u_core.u_sie._192_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._493_  (.A(\u_usb_host.u_core.status_rx_count_w[4] ),
    .B(net423),
    .X(\u_usb_host.u_core.u_sie._193_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._494_  (.A(\u_usb_host.u_core.status_rx_count_w[4] ),
    .B(net424),
    .Y(\u_usb_host.u_core.u_sie._194_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._495_  (.A(\u_usb_host.u_core.u_sie._193_ ),
    .B(\u_usb_host.u_core.u_sie._194_ ),
    .Y(\u_usb_host.u_core.u_sie._195_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._496_  (.A(\u_usb_host.u_core.u_sie._192_ ),
    .B(\u_usb_host.u_core.u_sie._195_ ),
    .Y(\u_usb_host.u_core.u_sie._196_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._497_  (.A(\u_usb_host.u_core.u_sie._192_ ),
    .B(\u_usb_host.u_core.u_sie._195_ ),
    .X(\u_usb_host.u_core.u_sie._197_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._498_  (.A1(net101),
    .A2(\u_usb_host.u_core.u_sie._196_ ),
    .A3(\u_usb_host.u_core.u_sie._197_ ),
    .B1(net106),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[4] ),
    .X(\u_usb_host.u_core.u_sie._010_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._499_  (.A(\u_usb_host.u_core.status_rx_count_w[5] ),
    .B(net424),
    .Y(\u_usb_host.u_core.u_sie._198_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_sie._500_  (.A(\u_usb_host.u_core.u_sie._194_ ),
    .B(\u_usb_host.u_core.u_sie._197_ ),
    .C(\u_usb_host.u_core.u_sie._198_ ),
    .Y(\u_usb_host.u_core.u_sie._199_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._501_  (.A1(\u_usb_host.u_core.u_sie._194_ ),
    .A2(\u_usb_host.u_core.u_sie._197_ ),
    .B1(\u_usb_host.u_core.u_sie._198_ ),
    .X(\u_usb_host.u_core.u_sie._200_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._502_  (.A1(net101),
    .A2(\u_usb_host.u_core.u_sie._199_ ),
    .A3(\u_usb_host.u_core.u_sie._200_ ),
    .B1(net106),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[5] ),
    .X(\u_usb_host.u_core.u_sie._011_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._503_  (.A(\u_usb_host.u_core.status_rx_count_w[6] ),
    .B(net423),
    .X(\u_usb_host.u_core.u_sie._201_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._504_  (.A(\u_usb_host.u_core.status_rx_count_w[6] ),
    .B(net423),
    .Y(\u_usb_host.u_core.u_sie._202_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._505_  (.A(\u_usb_host.u_core.u_sie._201_ ),
    .B(\u_usb_host.u_core.u_sie._202_ ),
    .Y(\u_usb_host.u_core.u_sie._203_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_sie._506_  (.A1(\u_usb_host.u_core.u_sie._101_ ),
    .A2(\u_usb_host.u_core.u_sie._121_ ),
    .B1(\u_usb_host.u_core.u_sie._197_ ),
    .B2(\u_usb_host.u_core.u_sie._198_ ),
    .X(\u_usb_host.u_core.u_sie._204_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie._507_  (.A(\u_usb_host.u_core.u_sie._203_ ),
    .B(\u_usb_host.u_core.u_sie._204_ ),
    .X(\u_usb_host.u_core.u_sie._205_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._508_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[6] ),
    .A2(net106),
    .B1(net101),
    .B2(\u_usb_host.u_core.u_sie._205_ ),
    .X(\u_usb_host.u_core.u_sie._012_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._509_  (.A1(\u_usb_host.u_core.u_sie._203_ ),
    .A2(\u_usb_host.u_core.u_sie._204_ ),
    .B1(\u_usb_host.u_core.u_sie._202_ ),
    .Y(\u_usb_host.u_core.u_sie._206_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._510_  (.A(\u_usb_host.u_core.status_rx_count_w[7] ),
    .B(net424),
    .Y(\u_usb_host.u_core.u_sie._207_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._511_  (.A(\u_usb_host.u_core.u_sie._206_ ),
    .B(\u_usb_host.u_core.u_sie._207_ ),
    .Y(\u_usb_host.u_core.u_sie._208_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._512_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[7] ),
    .A2(net106),
    .B1(net101),
    .B2(\u_usb_host.u_core.u_sie._208_ ),
    .X(\u_usb_host.u_core.u_sie._013_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._513_  (.A(\u_usb_host.u_core.u_sie._195_ ),
    .B(\u_usb_host.u_core.u_sie._198_ ),
    .C(\u_usb_host.u_core.u_sie._203_ ),
    .D(\u_usb_host.u_core.u_sie._207_ ),
    .X(\u_usb_host.u_core.u_sie._209_ ));
 sky130_fd_sc_hd__o2bb2a_1 \u_usb_host.u_core.u_sie._514_  (.A1_N(\u_usb_host.u_core.u_sie._102_ ),
    .A2_N(net424),
    .B1(\u_usb_host.u_core.u_sie._192_ ),
    .B2(\u_usb_host.u_core.u_sie._209_ ),
    .X(\u_usb_host.u_core.u_sie._210_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._515_  (.A(\u_usb_host.u_core.status_rx_count_w[8] ),
    .B(net423),
    .X(\u_usb_host.u_core.u_sie._211_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._516_  (.A(\u_usb_host.u_core.status_rx_count_w[8] ),
    .B(net423),
    .Y(\u_usb_host.u_core.u_sie._212_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._517_  (.A(\u_usb_host.u_core.u_sie._211_ ),
    .B(\u_usb_host.u_core.u_sie._212_ ),
    .Y(\u_usb_host.u_core.u_sie._213_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._518_  (.A(\u_usb_host.u_core.u_sie._210_ ),
    .B(\u_usb_host.u_core.u_sie._213_ ),
    .Y(\u_usb_host.u_core.u_sie._214_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._519_  (.A(\u_usb_host.u_core.u_sie._210_ ),
    .B(\u_usb_host.u_core.u_sie._213_ ),
    .X(\u_usb_host.u_core.u_sie._215_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._520_  (.A1(net101),
    .A2(\u_usb_host.u_core.u_sie._214_ ),
    .A3(\u_usb_host.u_core.u_sie._215_ ),
    .B1(net106),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[8] ),
    .X(\u_usb_host.u_core.u_sie._014_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._521_  (.A(\u_usb_host.u_core.status_rx_count_w[9] ),
    .B(net423),
    .Y(\u_usb_host.u_core.u_sie._216_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._522_  (.A1(\u_usb_host.u_core.u_sie._212_ ),
    .A2(\u_usb_host.u_core.u_sie._215_ ),
    .B1(\u_usb_host.u_core.u_sie._216_ ),
    .X(\u_usb_host.u_core.u_sie._217_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_sie._523_  (.A(\u_usb_host.u_core.u_sie._212_ ),
    .B(\u_usb_host.u_core.u_sie._215_ ),
    .C(\u_usb_host.u_core.u_sie._216_ ),
    .Y(\u_usb_host.u_core.u_sie._218_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._524_  (.A1(net101),
    .A2(\u_usb_host.u_core.u_sie._217_ ),
    .A3(\u_usb_host.u_core.u_sie._218_ ),
    .B1(net106),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[9] ),
    .X(\u_usb_host.u_core.u_sie._015_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._525_  (.A(\u_usb_host.u_core.status_rx_count_w[10] ),
    .B(net423),
    .X(\u_usb_host.u_core.u_sie._219_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._526_  (.A(\u_usb_host.u_core.status_rx_count_w[10] ),
    .B(net423),
    .Y(\u_usb_host.u_core.u_sie._220_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._527_  (.A(\u_usb_host.u_core.u_sie._219_ ),
    .B(\u_usb_host.u_core.u_sie._220_ ),
    .Y(\u_usb_host.u_core.u_sie._221_ ));
 sky130_fd_sc_hd__o22a_1 \u_usb_host.u_core.u_sie._528_  (.A1(\u_usb_host.u_core.u_sie._099_ ),
    .A2(\u_usb_host.u_core.u_sie._121_ ),
    .B1(\u_usb_host.u_core.u_sie._215_ ),
    .B2(\u_usb_host.u_core.u_sie._216_ ),
    .X(\u_usb_host.u_core.u_sie._222_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie._529_  (.A(\u_usb_host.u_core.u_sie._221_ ),
    .B(\u_usb_host.u_core.u_sie._222_ ),
    .X(\u_usb_host.u_core.u_sie._223_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._530_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[10] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._223_ ),
    .X(\u_usb_host.u_core.u_sie._001_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._531_  (.A1(\u_usb_host.u_core.u_sie._221_ ),
    .A2(\u_usb_host.u_core.u_sie._222_ ),
    .B1(\u_usb_host.u_core.u_sie._220_ ),
    .Y(\u_usb_host.u_core.u_sie._224_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._532_  (.A(\u_usb_host.u_core.status_rx_count_w[11] ),
    .B(net423),
    .Y(\u_usb_host.u_core.u_sie._225_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._533_  (.A(\u_usb_host.u_core.u_sie._224_ ),
    .B(\u_usb_host.u_core.u_sie._225_ ),
    .Y(\u_usb_host.u_core.u_sie._226_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._534_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[11] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._226_ ),
    .X(\u_usb_host.u_core.u_sie._002_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._535_  (.A(\u_usb_host.u_core.u_sie._213_ ),
    .B(\u_usb_host.u_core.u_sie._216_ ),
    .C(\u_usb_host.u_core.u_sie._221_ ),
    .D(\u_usb_host.u_core.u_sie._225_ ),
    .X(\u_usb_host.u_core.u_sie._227_ ));
 sky130_fd_sc_hd__o2bb2a_1 \u_usb_host.u_core.u_sie._536_  (.A1_N(\u_usb_host.u_core.u_sie._100_ ),
    .A2_N(net423),
    .B1(\u_usb_host.u_core.u_sie._210_ ),
    .B2(\u_usb_host.u_core.u_sie._227_ ),
    .X(\u_usb_host.u_core.u_sie._228_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._537_  (.A(\u_usb_host.u_core.status_rx_count_w[12] ),
    .B(net422),
    .X(\u_usb_host.u_core.u_sie._229_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._538_  (.A(\u_usb_host.u_core.status_rx_count_w[12] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._230_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._539_  (.A(\u_usb_host.u_core.u_sie._229_ ),
    .B(\u_usb_host.u_core.u_sie._230_ ),
    .Y(\u_usb_host.u_core.u_sie._231_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie._540_  (.A(\u_usb_host.u_core.u_sie._228_ ),
    .B(\u_usb_host.u_core.u_sie._231_ ),
    .X(\u_usb_host.u_core.u_sie._232_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._541_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[12] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._232_ ),
    .X(\u_usb_host.u_core.u_sie._003_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._542_  (.A1(\u_usb_host.u_core.u_sie._228_ ),
    .A2(\u_usb_host.u_core.u_sie._231_ ),
    .B1(\u_usb_host.u_core.u_sie._230_ ),
    .Y(\u_usb_host.u_core.u_sie._233_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._543_  (.A(\u_usb_host.u_core.status_rx_count_w[13] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._234_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._544_  (.A(\u_usb_host.u_core.u_sie._233_ ),
    .B(\u_usb_host.u_core.u_sie._234_ ),
    .Y(\u_usb_host.u_core.u_sie._235_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._545_  (.A1(\u_usb_host.u_core.u_sie.data_len_i[13] ),
    .A2(net105),
    .B1(net100),
    .B2(\u_usb_host.u_core.u_sie._235_ ),
    .X(\u_usb_host.u_core.u_sie._004_ ));
 sky130_fd_sc_hd__o32a_1 \u_usb_host.u_core.u_sie._546_  (.A1(\u_usb_host.u_core.u_sie._228_ ),
    .A2(\u_usb_host.u_core.u_sie._231_ ),
    .A3(\u_usb_host.u_core.u_sie._234_ ),
    .B1(\u_usb_host.u_core.u_sie._121_ ),
    .B2(\u_usb_host.u_core.u_sie._098_ ),
    .X(\u_usb_host.u_core.u_sie._236_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._547_  (.A(\u_usb_host.u_core.status_rx_count_w[14] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._237_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._548_  (.A(\u_usb_host.u_core.u_sie._237_ ),
    .Y(\u_usb_host.u_core.u_sie._238_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._549_  (.A(\u_usb_host.u_core.status_rx_count_w[14] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._239_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_core.u_sie._550_  (.A(\u_usb_host.u_core.u_sie._236_ ),
    .B(\u_usb_host.u_core.u_sie._238_ ),
    .C(\u_usb_host.u_core.u_sie._239_ ),
    .X(\u_usb_host.u_core.u_sie._240_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._551_  (.A1(\u_usb_host.u_core.u_sie._238_ ),
    .A2(\u_usb_host.u_core.u_sie._239_ ),
    .B1(\u_usb_host.u_core.u_sie._236_ ),
    .Y(\u_usb_host.u_core.u_sie._241_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._552_  (.A1(net100),
    .A2(\u_usb_host.u_core.u_sie._240_ ),
    .A3(\u_usb_host.u_core.u_sie._241_ ),
    .B1(net105),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[14] ),
    .X(\u_usb_host.u_core.u_sie._005_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie._553_  (.A(\u_usb_host.u_core.status_rx_count_w[15] ),
    .B(net422),
    .Y(\u_usb_host.u_core.u_sie._242_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._554_  (.A1(\u_usb_host.u_core.u_sie._237_ ),
    .A2(\u_usb_host.u_core.u_sie._240_ ),
    .B1(\u_usb_host.u_core.u_sie._242_ ),
    .X(\u_usb_host.u_core.u_sie._243_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_core.u_sie._555_  (.A(\u_usb_host.u_core.u_sie._237_ ),
    .B(\u_usb_host.u_core.u_sie._240_ ),
    .C(\u_usb_host.u_core.u_sie._242_ ),
    .Y(\u_usb_host.u_core.u_sie._244_ ));
 sky130_fd_sc_hd__a32o_1 \u_usb_host.u_core.u_sie._556_  (.A1(net100),
    .A2(\u_usb_host.u_core.u_sie._243_ ),
    .A3(\u_usb_host.u_core.u_sie._244_ ),
    .B1(net105),
    .B2(\u_usb_host.u_core.u_sie.data_len_i[15] ),
    .X(\u_usb_host.u_core.u_sie._006_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_core.u_sie._557_  (.A_N(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ),
    .B(\u_usb_host.u_core.u_sie._169_ ),
    .X(\u_usb_host.u_core.u_sie._033_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._558_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._245_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._559_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ),
    .B1(\u_usb_host.u_core.u_sie._245_ ),
    .Y(\u_usb_host.u_core.u_sie._034_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._560_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ),
    .B1(\u_usb_host.u_core.u_sie.last_tx_time_q[2] ),
    .X(\u_usb_host.u_core.u_sie._246_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_core.u_sie._561_  (.A_N(\u_usb_host.u_core.u_sie._124_ ),
    .B(\u_usb_host.u_core.u_sie._169_ ),
    .C(\u_usb_host.u_core.u_sie._246_ ),
    .X(\u_usb_host.u_core.u_sie._035_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._562_  (.A(\u_usb_host.u_core.u_sie.last_tx_time_q[3] ),
    .B(\u_usb_host.u_core.u_sie._124_ ),
    .X(\u_usb_host.u_core.u_sie._247_ ));
 sky130_fd_sc_hd__and3b_1 \u_usb_host.u_core.u_sie._563_  (.A_N(\u_usb_host.u_core.u_sie._125_ ),
    .B(\u_usb_host.u_core.u_sie._169_ ),
    .C(\u_usb_host.u_core.u_sie._247_ ),
    .X(\u_usb_host.u_core.u_sie._036_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._564_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[4] ),
    .A2(\u_usb_host.u_core.u_sie._125_ ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._248_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._565_  (.A(\u_usb_host.u_core.u_sie._126_ ),
    .B(\u_usb_host.u_core.u_sie._248_ ),
    .Y(\u_usb_host.u_core.u_sie._037_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._566_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[5] ),
    .A2(\u_usb_host.u_core.u_sie._126_ ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._249_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._567_  (.A(\u_usb_host.u_core.u_sie._127_ ),
    .B(\u_usb_host.u_core.u_sie._249_ ),
    .Y(\u_usb_host.u_core.u_sie._038_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._568_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[6] ),
    .A2(\u_usb_host.u_core.u_sie._127_ ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._250_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._569_  (.A(\u_usb_host.u_core.u_sie._128_ ),
    .B(\u_usb_host.u_core.u_sie._250_ ),
    .Y(\u_usb_host.u_core.u_sie._039_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._570_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[7] ),
    .A2(\u_usb_host.u_core.u_sie._128_ ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._251_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._571_  (.A(\u_usb_host.u_core.u_sie._129_ ),
    .B(\u_usb_host.u_core.u_sie._251_ ),
    .Y(\u_usb_host.u_core.u_sie._040_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._572_  (.A1(\u_usb_host.u_core.u_sie.last_tx_time_q[8] ),
    .A2(\u_usb_host.u_core.u_sie._129_ ),
    .B1(\u_usb_host.u_core.u_sie._169_ ),
    .Y(\u_usb_host.u_core.u_sie._252_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._573_  (.A(\u_usb_host.u_core.u_sie._130_ ),
    .B(\u_usb_host.u_core.u_sie._252_ ),
    .Y(\u_usb_host.u_core.u_sie._041_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._574_  (.A(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ),
    .B(net582),
    .Y(\u_usb_host.u_core.u_sie._059_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._575_  (.A1(\u_usb_host.u_core.u_sie.tx_ifs_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ),
    .B1(net582),
    .Y(\u_usb_host.u_core.u_sie._253_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._576_  (.A1(\u_usb_host.u_core.u_sie.tx_ifs_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ),
    .B1(\u_usb_host.u_core.u_sie._253_ ),
    .Y(\u_usb_host.u_core.u_sie._060_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._577_  (.A1(\u_usb_host.u_core.u_sie.tx_ifs_q[1] ),
    .A2(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ),
    .B1(\u_usb_host.u_core.u_sie.tx_ifs_q[2] ),
    .Y(\u_usb_host.u_core.u_sie._254_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._578_  (.A1(\u_usb_host.u_core.u_sie._093_ ),
    .A2(\u_usb_host.u_core.u_sie._254_ ),
    .B1(net582),
    .Y(\u_usb_host.u_core.u_sie._061_ ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._579_  (.A1(\u_usb_host.u_core.u_sie.tx_ifs_q[3] ),
    .A2(\u_usb_host.u_core.u_sie._093_ ),
    .B1(net582),
    .Y(\u_usb_host.u_core.u_sie._255_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._580_  (.A(\u_usb_host.u_core.u_sie._094_ ),
    .B(\u_usb_host.u_core.u_sie._255_ ),
    .Y(\u_usb_host.u_core.u_sie._062_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._581_  (.A1(net425),
    .A2(\u_usb_host.u_core.fifo_tx_data_w[0] ),
    .B1(\u_usb_host.u_core.u_sie._097_ ),
    .X(\u_usb_host.u_core.u_sie._256_ ));
 sky130_fd_sc_hd__a221o_1 \u_usb_host.u_core.u_sie._582_  (.A1(\u_usb_host.u_core.u_sie.token_q[7] ),
    .A2(\u_usb_host.u_core.u_sie._107_ ),
    .B1(\u_usb_host.u_core.u_sie._139_ ),
    .B2(\u_usb_host.u_core.u_sie.token_q[15] ),
    .C1(\u_usb_host.u_core.u_sie._256_ ),
    .X(\u_usb_host.u_core.u_sie._257_ ));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_core.u_sie._583_  (.A1(\u_usb_host.u_core.u_sie.crc_sum_q[8] ),
    .A2(\u_usb_host.u_core.u_sie._091_ ),
    .B1(\u_usb_host.u_core.u_sie._116_ ),
    .B2(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .Y(\u_usb_host.u_core.u_sie._258_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._584_  (.A1(\u_usb_host.u_core.token_pid_w[0] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._257_ ),
    .C1(\u_usb_host.u_core.u_sie._258_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[0] ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._585_  (.A1(net425),
    .A2(\u_usb_host.u_core.u_sie._097_ ),
    .B1(\u_usb_host.u_core.u_sie._105_ ),
    .X(\u_usb_host.u_core.u_sie._259_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._586_  (.A1(\u_usb_host.u_core.fifo_tx_data_w[1] ),
    .A2(\u_usb_host.u_core.u_sie._147_ ),
    .B1(\u_usb_host.u_core.u_sie._259_ ),
    .X(\u_usb_host.u_core.u_sie._260_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._587_  (.A(\u_usb_host.u_core.u_sie.token_q[6] ),
    .B(\u_usb_host.u_core.u_sie._108_ ),
    .X(\u_usb_host.u_core.u_sie._261_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._588_  (.A1(\u_usb_host.u_core.u_sie.token_q[14] ),
    .A2(\u_usb_host.u_core.u_sie._139_ ),
    .B1(\u_usb_host.u_core.u_sie._260_ ),
    .B2(\u_usb_host.u_core.u_sie._261_ ),
    .X(\u_usb_host.u_core.u_sie._262_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._589_  (.A1(\u_usb_host.u_core.token_pid_w[1] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._262_ ),
    .C1(\u_usb_host.u_core.u_sie._292_ ),
    .X(\u_usb_host.u_core.u_sie._263_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._590_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[9] ),
    .B(\u_usb_host.u_core.u_sie._292_ ),
    .Y(\u_usb_host.u_core.u_sie._264_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_sie._591_  (.A1_N(\u_usb_host.u_core.u_sie.crc_sum_q[1] ),
    .A2_N(\u_usb_host.u_core.u_sie._116_ ),
    .B1(\u_usb_host.u_core.u_sie._263_ ),
    .B2(\u_usb_host.u_core.u_sie._264_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[1] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._592_  (.A1(\u_usb_host.u_core.u_sie.token_q[5] ),
    .A2(\u_usb_host.u_core.u_sie._107_ ),
    .B1(\u_usb_host.u_core.u_sie._147_ ),
    .B2(\u_usb_host.u_core.fifo_tx_data_w[2] ),
    .X(\u_usb_host.u_core.u_sie._265_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._593_  (.A0(\u_usb_host.u_core.u_sie._265_ ),
    .A1(\u_usb_host.u_core.u_sie.token_q[13] ),
    .S(\u_usb_host.u_core.u_sie._139_ ),
    .X(\u_usb_host.u_core.u_sie._266_ ));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_core.u_sie._594_  (.A1(\u_usb_host.u_core.u_sie.crc_sum_q[10] ),
    .A2(\u_usb_host.u_core.u_sie._091_ ),
    .B1(\u_usb_host.u_core.u_sie._116_ ),
    .B2(\u_usb_host.u_core.u_sie.crc_sum_q[2] ),
    .Y(\u_usb_host.u_core.u_sie._267_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._595_  (.A1(\u_usb_host.u_core.token_pid_w[2] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._266_ ),
    .C1(\u_usb_host.u_core.u_sie._267_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[2] ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_core.u_sie._596_  (.A1(net425),
    .A2(\u_usb_host.u_core.u_sie.send_data1_q ),
    .A3(\u_usb_host.u_core.u_sie._097_ ),
    .B1(\u_usb_host.u_core.u_sie._107_ ),
    .X(\u_usb_host.u_core.u_sie._268_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._597_  (.A1(\u_usb_host.u_core.fifo_tx_data_w[3] ),
    .A2(\u_usb_host.u_core.u_sie._147_ ),
    .B1(\u_usb_host.u_core.u_sie._268_ ),
    .X(\u_usb_host.u_core.u_sie._269_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._598_  (.A(\u_usb_host.u_core.u_sie.token_q[4] ),
    .B(\u_usb_host.u_core.u_sie._108_ ),
    .X(\u_usb_host.u_core.u_sie._270_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._599_  (.A1(\u_usb_host.u_core.u_sie.token_q[12] ),
    .A2(\u_usb_host.u_core.u_sie._139_ ),
    .B1(\u_usb_host.u_core.u_sie._269_ ),
    .B2(\u_usb_host.u_core.u_sie._270_ ),
    .X(\u_usb_host.u_core.u_sie._271_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._600_  (.A1(\u_usb_host.u_core.token_pid_w[3] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._271_ ),
    .C1(\u_usb_host.u_core.u_sie._292_ ),
    .X(\u_usb_host.u_core.u_sie._272_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._601_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[11] ),
    .B(\u_usb_host.u_core.u_sie._292_ ),
    .Y(\u_usb_host.u_core.u_sie._273_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_sie._602_  (.A1_N(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .A2_N(\u_usb_host.u_core.u_sie._116_ ),
    .B1(\u_usb_host.u_core.u_sie._272_ ),
    .B2(\u_usb_host.u_core.u_sie._273_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[3] ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._603_  (.A1(\u_usb_host.u_core.fifo_tx_data_w[4] ),
    .A2(\u_usb_host.u_core.u_sie._147_ ),
    .B1(\u_usb_host.u_core.u_sie._105_ ),
    .X(\u_usb_host.u_core.u_sie._274_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_core.u_sie._604_  (.A1(\u_usb_host.u_core.u_sie.token_q[3] ),
    .A2(\u_usb_host.u_core.u_sie._108_ ),
    .B1(\u_usb_host.u_core.u_sie._274_ ),
    .X(\u_usb_host.u_core.u_sie._275_ ));
 sky130_fd_sc_hd__a221oi_2 \u_usb_host.u_core.u_sie._605_  (.A1(\u_usb_host.u_core.token_pid_w[4] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._139_ ),
    .B2(\u_usb_host.u_core.u_sie.token_q[11] ),
    .C1(\u_usb_host.u_core.u_sie._275_ ),
    .Y(\u_usb_host.u_core.u_sie._276_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._606_  (.A0(\u_usb_host.u_core.u_sie.crc_sum_q[12] ),
    .A1(\u_usb_host.u_core.u_sie._276_ ),
    .S(\u_usb_host.u_core.u_sie._091_ ),
    .X(\u_usb_host.u_core.u_sie._277_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_core.u_sie._607_  (.A1(\u_usb_host.u_core.u_sie.crc_sum_q[4] ),
    .A2(\u_usb_host.u_core.u_sie._116_ ),
    .B1(\u_usb_host.u_core.u_sie._277_ ),
    .Y(\u_usb_host.u_core.u_sie.utmi_data_o[4] ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._608_  (.A1(\u_usb_host.u_core.u_sie.token_q[2] ),
    .A2(\u_usb_host.u_core.u_sie._107_ ),
    .B1(\u_usb_host.u_core.u_sie._147_ ),
    .B2(\u_usb_host.u_core.fifo_tx_data_w[5] ),
    .X(\u_usb_host.u_core.u_sie._278_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._609_  (.A0(\u_usb_host.u_core.u_sie._278_ ),
    .A1(\u_usb_host.u_core.u_sie.token_q[10] ),
    .S(\u_usb_host.u_core.u_sie._139_ ),
    .X(\u_usb_host.u_core.u_sie._279_ ));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_core.u_sie._610_  (.A1(\u_usb_host.u_core.u_sie.crc_sum_q[13] ),
    .A2(\u_usb_host.u_core.u_sie._091_ ),
    .B1(\u_usb_host.u_core.u_sie._116_ ),
    .B2(\u_usb_host.u_core.u_sie.crc_sum_q[5] ),
    .Y(\u_usb_host.u_core.u_sie._280_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._611_  (.A1(\u_usb_host.u_core.token_pid_w[5] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._279_ ),
    .C1(\u_usb_host.u_core.u_sie._280_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[5] ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._612_  (.A1(\u_usb_host.u_core.fifo_tx_data_w[6] ),
    .A2(\u_usb_host.u_core.u_sie._147_ ),
    .B1(\u_usb_host.u_core.u_sie._259_ ),
    .X(\u_usb_host.u_core.u_sie._281_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_core.u_sie._613_  (.A(\u_usb_host.u_core.u_sie.token_q[1] ),
    .B(\u_usb_host.u_core.u_sie._108_ ),
    .X(\u_usb_host.u_core.u_sie._282_ ));
 sky130_fd_sc_hd__a22o_1 \u_usb_host.u_core.u_sie._614_  (.A1(\u_usb_host.u_core.u_sie.token_q[9] ),
    .A2(\u_usb_host.u_core.u_sie._139_ ),
    .B1(\u_usb_host.u_core.u_sie._281_ ),
    .B2(\u_usb_host.u_core.u_sie._282_ ),
    .X(\u_usb_host.u_core.u_sie._283_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._615_  (.A1(\u_usb_host.u_core.token_pid_w[6] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._283_ ),
    .C1(\u_usb_host.u_core.u_sie._292_ ),
    .X(\u_usb_host.u_core.u_sie._284_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_core.u_sie._616_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[14] ),
    .B(\u_usb_host.u_core.u_sie._292_ ),
    .Y(\u_usb_host.u_core.u_sie._285_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._617_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[6] ),
    .B(\u_usb_host.u_core.u_sie._116_ ),
    .Y(\u_usb_host.u_core.u_sie._286_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_core.u_sie._618_  (.A1(\u_usb_host.u_core.u_sie._284_ ),
    .A2(\u_usb_host.u_core.u_sie._285_ ),
    .B1(\u_usb_host.u_core.u_sie._286_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[6] ));
 sky130_fd_sc_hd__a21oi_1 \u_usb_host.u_core.u_sie._619_  (.A1(\u_usb_host.u_core.fifo_tx_data_w[7] ),
    .A2(\u_usb_host.u_core.u_sie._147_ ),
    .B1(\u_usb_host.u_core.u_sie._259_ ),
    .Y(\u_usb_host.u_core.u_sie._287_ ));
 sky130_fd_sc_hd__a2bb2o_1 \u_usb_host.u_core.u_sie._620_  (.A1_N(\u_usb_host.u_core.u_sie._268_ ),
    .A2_N(\u_usb_host.u_core.u_sie._287_ ),
    .B1(\u_usb_host.u_core.u_sie.token_q[0] ),
    .B2(\u_usb_host.u_core.u_sie._107_ ),
    .X(\u_usb_host.u_core.u_sie._288_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._621_  (.A0(\u_usb_host.u_core.u_sie._288_ ),
    .A1(\u_usb_host.u_core.u_sie.token_q[8] ),
    .S(\u_usb_host.u_core.u_sie._139_ ),
    .X(\u_usb_host.u_core.u_sie._289_ ));
 sky130_fd_sc_hd__o22ai_1 \u_usb_host.u_core.u_sie._622_  (.A1(\u_usb_host.u_core.u_sie.crc_sum_q[15] ),
    .A2(\u_usb_host.u_core.u_sie._091_ ),
    .B1(\u_usb_host.u_core.u_sie._116_ ),
    .B2(\u_usb_host.u_core.u_sie.crc_sum_q[7] ),
    .Y(\u_usb_host.u_core.u_sie._290_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_core.u_sie._623_  (.A1(\u_usb_host.u_core.token_pid_w[7] ),
    .A2(\u_usb_host.u_core.u_sie._117_ ),
    .B1(\u_usb_host.u_core.u_sie._289_ ),
    .C1(\u_usb_host.u_core.u_sie._290_ ),
    .X(\u_usb_host.u_core.u_sie.utmi_data_o[7] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._624_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[0] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[0] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[0] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._625_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[1] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[1] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[1] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._626_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[2] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[2] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[2] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._627_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[3] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[3] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[3] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._628_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[4] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[4] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[4] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._629_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[5] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[5] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[5] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._630_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[6] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[6] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[6] ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_core.u_sie._631_  (.A0(\u_usb_host.u_core.u_sie.data_buffer_q[7] ),
    .A1(\u_usb_host.u_core.fifo_tx_data_w[7] ),
    .S(net183),
    .X(\u_usb_host.u_core.u_sie.crc_data_in_w[7] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._632_  (.A(\u_usb_host.u_core.u_sie._292_ ),
    .B(\u_usb_host.u_core.u_sie._123_ ),
    .Y(\u_usb_host.u_core.u_sie._073_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_core.u_sie._633_  (.A(\u_usb_host.u_core.u_sie.data_valid_q[1] ),
    .B(\u_usb_host.u_core.u_sie.shift_en_w ),
    .X(\u_usb_host.u_core.u_sie._032_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_core.u_sie._634_  (.A(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .B(net183),
    .Y(\u_usb_host.u_core.u_sie._052_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_core.u_sie._635_  (.A(\u_usb_host.u_core.u_sie._083_ ),
    .B(\u_usb_host.u_core.u_sie.crc_byte_w ),
    .C(net114),
    .D(\u_usb_host.u_core.u_sie._123_ ),
    .X(\u_usb_host.u_core.u_sie._291_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_core.u_sie._636_  (.A(\u_usb_host.u_core.u_sie._291_ ),
    .Y(\u_usb_host.u_core.fifo_rx_push_w ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._637_  (.CLK(clknet_leaf_16_usb_clk),
    .D(\u_usb_host.u_core.u_sie._032_ ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_ready_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._638_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_ep_w[0] ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.u_sie.token_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._639_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_ep_w[1] ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.u_sie.token_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._640_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_ep_w[2] ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.u_sie.token_q[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._641_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_ep_w[3] ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.u_sie.token_q[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._642_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[0] ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.u_sie.token_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._643_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[1] ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.u_sie.token_q[10] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._644_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[2] ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.u_sie.token_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._645_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[3] ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.u_sie.token_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._646_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[4] ),
    .RESET_B(net376),
    .Q(\u_usb_host.u_core.u_sie.token_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._647_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[5] ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.u_sie.token_q[14] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._648_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._310_ ),
    .D(\u_usb_host.u_core.token_dev_w[6] ),
    .RESET_B(net375),
    .Q(\u_usb_host.u_core.u_sie.token_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._649_  (.CLK(\u_usb_host.u_core.u_sie._298_ ),
    .D(net688),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.u_sie.send_data1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._650_  (.CLK(\u_usb_host.u_core.u_sie._299_ ),
    .D(net525),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.u_sie.send_sof_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._651_  (.CLK(\u_usb_host.u_core.u_sie._300_ ),
    .D(\u_usb_host.u_core.u_sie._079_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.u_sie.send_ack_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._652_  (.CLK(\u_usb_host.u_core.u_sie._309_ ),
    .D(\u_usb_host.u_core.u_sie._043_ ),
    .RESET_B(net403),
    .Q(\u_usb_host.u_core.status_crc_err_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._653_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._311_ ),
    .D(\u_usb_host.u_core.u_sie._054_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.token_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._654_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._311_ ),
    .D(\u_usb_host.u_core.u_sie._055_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.token_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._655_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._311_ ),
    .D(\u_usb_host.u_core.u_sie._056_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_sie.token_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._656_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._311_ ),
    .D(\u_usb_host.u_core.u_sie._057_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.token_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._657_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._311_ ),
    .D(\u_usb_host.u_core.u_sie._058_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.token_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._658_  (.CLK(\u_usb_host.u_core.u_sie._293_ ),
    .D(\u_usb_host.u_core.u_sie._063_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.wait_eop_q ));
 sky130_fd_sc_hd__dfstp_2 \u_usb_host.u_core.u_sie._659_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._016_ ),
    .SET_B(net411),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[0] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._660_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._023_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[1] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._661_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._024_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[2] ));
 sky130_fd_sc_hd__dfstp_2 \u_usb_host.u_core.u_sie._662_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._025_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[3] ));
 sky130_fd_sc_hd__dfstp_2 \u_usb_host.u_core.u_sie._663_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._026_ ),
    .SET_B(net402),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[4] ));
 sky130_fd_sc_hd__dfstp_2 \u_usb_host.u_core.u_sie._664_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._027_ ),
    .SET_B(net402),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[5] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._665_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._028_ ),
    .SET_B(net402),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[6] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._666_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._029_ ),
    .SET_B(net402),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[7] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._667_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._030_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[8] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._668_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._031_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[9] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._669_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._017_ ),
    .SET_B(net405),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[10] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._670_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._018_ ),
    .SET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[11] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._671_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._019_ ),
    .SET_B(net402),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[12] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._672_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._020_ ),
    .SET_B(net401),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[13] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._673_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._021_ ),
    .SET_B(net401),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[14] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_core.u_sie._674_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._312_ ),
    .D(\u_usb_host.u_core.u_sie._022_ ),
    .SET_B(net411),
    .Q(\u_usb_host.u_core.u_sie.crc_sum_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._675_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._294_ ),
    .D(\u_usb_host.u_core.u_sie._059_ ),
    .RESET_B(net409),
    .Q(\u_usb_host.u_core.u_sie.tx_ifs_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._676_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._294_ ),
    .D(\u_usb_host.u_core.u_sie._060_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.tx_ifs_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._677_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._294_ ),
    .D(\u_usb_host.u_core.u_sie._061_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.tx_ifs_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._678_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._294_ ),
    .D(\u_usb_host.u_core.u_sie._062_ ),
    .RESET_B(net409),
    .Q(\u_usb_host.u_core.u_sie.tx_ifs_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._679_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._033_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._680_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._034_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._681_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._035_ ),
    .RESET_B(net400),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._682_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._036_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._683_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._037_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._684_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._038_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._685_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._039_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._686_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._040_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._687_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._295_ ),
    .D(\u_usb_host.u_core.u_sie._041_ ),
    .RESET_B(net399),
    .Q(\u_usb_host.u_core.u_sie.last_tx_time_q[8] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._688_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._000_ ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.status_rx_count_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._689_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._007_ ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.status_rx_count_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._690_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._008_ ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.status_rx_count_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._691_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._009_ ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.status_rx_count_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._692_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._010_ ),
    .RESET_B(net393),
    .Q(\u_usb_host.u_core.status_rx_count_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._693_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._011_ ),
    .RESET_B(net394),
    .Q(\u_usb_host.u_core.status_rx_count_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._694_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._012_ ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.status_rx_count_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._695_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._013_ ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.status_rx_count_w[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._696_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._014_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._697_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._015_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._698_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._001_ ),
    .RESET_B(net385),
    .Q(\u_usb_host.u_core.status_rx_count_w[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._699_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._002_ ),
    .RESET_B(net385),
    .Q(\u_usb_host.u_core.status_rx_count_w[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._700_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._003_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[12] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._701_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._004_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._702_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._005_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._703_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._296_ ),
    .D(\u_usb_host.u_core.u_sie._006_ ),
    .RESET_B(net384),
    .Q(\u_usb_host.u_core.status_rx_count_w[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._704_  (.CLK(\u_usb_host.u_core.u_sie._297_ ),
    .D(net684),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.u_sie.in_transfer_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._705_  (.CLK(\u_usb_host.u_core.u_sie._301_ ),
    .D(\u_usb_host.u_core.u_sie._064_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.u_sie.wait_resp_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._706_  (.CLK(\u_usb_host.u_core.u_sie._302_ ),
    .D(\u_usb_host.u_core.u_sie._292_ ),
    .RESET_B(net405),
    .Q(\u_usb_host.u_core.status_tx_done_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._707_  (.CLK(\u_usb_host.u_core.u_sie._303_ ),
    .D(\u_usb_host.u_core.u_sie._052_ ),
    .RESET_B(net405),
    .Q(\u_usb_host.u_core.status_rx_done_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._708_  (.CLK(\u_usb_host.u_core.u_sie._304_ ),
    .D(\u_usb_host.u_core.u_sie._053_ ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.status_timeout_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._709_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._044_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.status_response_w[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._710_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._045_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.status_response_w[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._711_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._046_ ),
    .RESET_B(net398),
    .Q(\u_usb_host.u_core.status_response_w[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._712_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._047_ ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.status_response_w[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._713_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._048_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.status_response_w[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._714_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._049_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.status_response_w[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._715_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._050_ ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.status_response_w[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._716_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._305_ ),
    .D(\u_usb_host.u_core.u_sie._051_ ),
    .RESET_B(net396),
    .Q(\u_usb_host.u_core.status_response_w[7] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._717_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net637),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[0] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._718_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net651),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._719_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net639),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._720_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net653),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._721_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net652),
    .RESET_B(net411),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[4] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._722_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net650),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._723_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net672),
    .RESET_B(net411),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[6] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._724_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net665),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._725_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net667),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[8] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._726_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net634),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[9] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._727_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net638),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[10] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._728_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net633),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[11] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._729_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net642),
    .RESET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[12] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._730_  (.CLK(\clknet_2_3__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net635),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[13] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._731_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net649),
    .RESET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[14] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._732_  (.CLK(\clknet_2_1__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net636),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[15] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._733_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net663),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[16] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._734_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net666),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[17] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._735_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net661),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[18] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._736_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net664),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[19] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._737_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net654),
    .RESET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[20] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._738_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net670),
    .RESET_B(net412),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[21] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._739_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net669),
    .RESET_B(net410),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[22] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._740_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net662),
    .RESET_B(net413),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[23] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._741_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[24] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._742_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net622),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[25] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._743_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net616),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[26] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._744_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net611),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[27] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._745_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net620),
    .RESET_B(net405),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[28] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._746_  (.CLK(\clknet_2_2__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net621),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[29] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._747_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net624),
    .RESET_B(net405),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[30] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._748_  (.CLK(\clknet_2_0__leaf_u_usb_host.u_core.u_sie._306_ ),
    .D(net615),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.data_buffer_q[31] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._749_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._307_ ),
    .D(net660),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_valid_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._750_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._307_ ),
    .D(net631),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_valid_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._751_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._307_ ),
    .D(\u_usb_host.u_core.u_sie._065_ ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.data_valid_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._752_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_core.u_sie._308_ ),
    .D(net641),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.crc_byte_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._753_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_core.u_sie._308_ ),
    .D(\u_usb_host.u_core.u_sie._080_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.data_crc_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._754_  (.CLK(clknet_leaf_17_usb_clk),
    .D(\u_usb_host.u_core.u_sie.next_state_r[0] ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._755_  (.CLK(clknet_leaf_18_usb_clk),
    .D(\u_usb_host.u_core.u_sie.next_state_r[1] ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.state_q[1] ));
 sky130_fd_sc_hd__dfrtp_4 \u_usb_host.u_core.u_sie._756_  (.CLK(clknet_leaf_18_usb_clk),
    .D(\u_usb_host.u_core.u_sie.next_state_r[2] ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.state_q[2] ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_core.u_sie._757_  (.CLK(clknet_leaf_18_usb_clk),
    .D(\u_usb_host.u_core.u_sie.next_state_r[3] ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.state_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._758_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.u_sie.utmi_linestate_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._759_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.u_sie.utmi_linestate_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._760_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_core.u_sie.se0_detect_w ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.u_sie.se0_detect_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._761_  (.CLK(clknet_leaf_19_usb_clk),
    .D(\u_usb_host.u_core.u_sie._042_ ),
    .RESET_B(net397),
    .Q(\u_usb_host.u_core.transfer_ack_w ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._762_  (.CLK(clknet_leaf_17_usb_clk),
    .D(net675),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.rx_active_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._763_  (.CLK(clknet_leaf_15_usb_clk),
    .D(net676),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.rx_active_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._764_  (.CLK(clknet_leaf_15_usb_clk),
    .D(\u_usb_host.u_core.u_sie.rx_active_q[3] ),
    .RESET_B(net404),
    .Q(\u_usb_host.u_core.u_sie.rx_active_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_core.u_sie._765_  (.CLK(clknet_leaf_15_usb_clk),
    .D(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.rx_active_q[3] ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._766_  (.CLK(clknet_leaf_15_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._066_ ),
    .GCLK(\u_usb_host.u_core.u_sie._293_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._767_  (.CLK(clknet_leaf_15_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._067_ ),
    .GCLK(\u_usb_host.u_core.u_sie._294_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._768_  (.CLK(clknet_leaf_20_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._068_ ),
    .GCLK(\u_usb_host.u_core.u_sie._295_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._769_  (.CLK(clknet_leaf_13_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._069_ ),
    .GCLK(\u_usb_host.u_core.u_sie._296_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._770_  (.CLK(clknet_leaf_19_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._070_ ),
    .GCLK(\u_usb_host.u_core.u_sie._297_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._771_  (.CLK(clknet_leaf_19_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._070_ ),
    .GCLK(\u_usb_host.u_core.u_sie._298_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._772_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._070_ ),
    .GCLK(\u_usb_host.u_core.u_sie._299_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._773_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._070_ ),
    .GCLK(\u_usb_host.u_core.u_sie._300_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._774_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._071_ ),
    .GCLK(\u_usb_host.u_core.u_sie._301_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._775_  (.CLK(clknet_leaf_17_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._072_ ),
    .GCLK(\u_usb_host.u_core.u_sie._302_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._776_  (.CLK(clknet_leaf_17_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._073_ ),
    .GCLK(\u_usb_host.u_core.u_sie._303_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._777_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._074_ ),
    .GCLK(\u_usb_host.u_core.u_sie._304_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._778_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._075_ ),
    .GCLK(\u_usb_host.u_core.u_sie._305_ ));
 sky130_fd_sc_hd__dlclkp_4 \u_usb_host.u_core.u_sie._779_  (.CLK(clknet_leaf_16_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie.shift_en_w ),
    .GCLK(\u_usb_host.u_core.u_sie._306_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._780_  (.CLK(clknet_leaf_15_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie.shift_en_w ),
    .GCLK(\u_usb_host.u_core.u_sie._307_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._781_  (.CLK(clknet_leaf_15_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie.shift_en_w ),
    .GCLK(\u_usb_host.u_core.u_sie._308_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_core.u_sie._782_  (.CLK(clknet_leaf_18_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._076_ ),
    .GCLK(\u_usb_host.u_core.u_sie._309_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._783_  (.CLK(clknet_leaf_19_usb_clk),
    .GATE(net113),
    .GCLK(\u_usb_host.u_core.u_sie._310_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._784_  (.CLK(clknet_leaf_21_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._077_ ),
    .GCLK(\u_usb_host.u_core.u_sie._311_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_core.u_sie._785_  (.CLK(clknet_leaf_17_usb_clk),
    .GATE(\u_usb_host.u_core.u_sie._078_ ),
    .GCLK(\u_usb_host.u_core.u_sie._312_ ));
 sky130_fd_sc_hd__clkbuf_2 \u_usb_host.u_core.u_sie._791_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[0] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[0] ));
 sky130_fd_sc_hd__clkbuf_4 \u_usb_host.u_core.u_sie._792_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[1] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[1] ));
 sky130_fd_sc_hd__clkbuf_2 \u_usb_host.u_core.u_sie._793_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[2] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[2] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._794_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[3] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[3] ));
 sky130_fd_sc_hd__clkbuf_2 \u_usb_host.u_core.u_sie._795_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[4] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[4] ));
 sky130_fd_sc_hd__buf_2 \u_usb_host.u_core.u_sie._796_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[5] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[5] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._797_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[6] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[6] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie._798_  (.A(\u_usb_host.u_core.u_sie.data_buffer_q[7] ),
    .X(\u_usb_host.u_core.fifo_rx_data_w[7] ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc16._29_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[2] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[1] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._00_ ));
 sky130_fd_sc_hd__xnor2_2 \u_usb_host.u_core.u_sie.u_crc16._30_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[4] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._00_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._01_ ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc16._31_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[1] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[0] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._02_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._32_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[5] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._02_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._03_ ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc16._33_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[2] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[3] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._04_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._34_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[4] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[6] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._05_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._35_  (.A(\u_usb_host.u_core.u_sie.u_crc16._04_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._05_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._06_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._36_  (.A(\u_usb_host.u_core.u_sie.u_crc16._03_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._06_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._07_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._37_  (.A(\u_usb_host.u_core.u_sie.u_crc16._01_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._07_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._08_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._38_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[5] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._09_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._39_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[7] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._09_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._10_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._40_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[7] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[6] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._11_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._41_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._11_ ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._12_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._42_  (.A(\u_usb_host.u_core.u_sie.u_crc16._10_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._12_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._13_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._43_  (.A(\u_usb_host.u_core.u_sie.u_crc16._08_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._13_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[15] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._44_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[6] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[5] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._14_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._45_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._15_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._46_  (.A(\u_usb_host.u_core.u_sie.u_crc16._14_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._15_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._16_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._47_  (.A(\u_usb_host.u_core.u_sie.u_crc16._01_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._16_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._17_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._48_  (.A(\u_usb_host.u_core.u_sie.u_crc16._07_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._17_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[14] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._49_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[6] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[7] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._18_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._50_  (.A(\u_usb_host.u_core.u_sie.u_crc16._11_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._18_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[13] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._51_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[5] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[6] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._19_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._52_  (.A(\u_usb_host.u_core.u_sie.u_crc16._14_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._19_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[12] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._53_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[5] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[4] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._20_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._54_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[4] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[5] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._21_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._55_  (.A(\u_usb_host.u_core.u_sie.u_crc16._20_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._21_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[11] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._56_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[4] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._22_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._57_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[3] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[4] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._23_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._58_  (.A(\u_usb_host.u_core.u_sie.u_crc16._22_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._23_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[10] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._59_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[3] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[2] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._24_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._60_  (.A(\u_usb_host.u_core.u_sie.u_crc16._04_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._24_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[9] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._61_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[1] ),
    .B(\u_usb_host.u_core.u_sie.crc_data_in_w[2] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._25_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._62_  (.A(\u_usb_host.u_core.u_sie.u_crc16._00_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._25_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[8] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._63_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[1] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[15] ),
    .X(\u_usb_host.u_core.u_sie.u_crc16._26_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._64_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._26_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._27_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._65_  (.A(\u_usb_host.u_core.u_sie.u_crc16._02_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._27_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[7] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._66_  (.A(\u_usb_host.u_core.u_sie.crc_data_in_w[0] ),
    .B(\u_usb_host.u_core.u_sie.crc_sum_q[14] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc16._28_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc16._67_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[0] ),
    .B(\u_usb_host.u_core.u_sie.u_crc16._28_ ),
    .Y(\u_usb_host.u_core.u_sie.crc_out_w[6] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc16._68_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[8] ),
    .B(\u_usb_host.u_core.u_sie.crc_out_w[15] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[0] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie.u_crc16._69_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[9] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[1] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie.u_crc16._70_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[10] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[2] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie.u_crc16._71_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[11] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[3] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie.u_crc16._72_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[12] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[4] ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_core.u_sie.u_crc16._73_  (.A(\u_usb_host.u_core.u_sie.crc_sum_q[13] ),
    .X(\u_usb_host.u_core.u_sie.crc_out_w[5] ));
 sky130_fd_sc_hd__xnor2_2 \u_usb_host.u_core.u_sie.u_crc5._29_  (.A(\u_usb_host.u_core.u_sie.token_q[14] ),
    .B(\u_usb_host.u_core.u_sie.token_q[15] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._00_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._30_  (.A(\u_usb_host.u_core.u_sie.token_q[5] ),
    .B(net556),
    .X(\u_usb_host.u_core.u_sie.u_crc5._01_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._30__556  (.HI(net556));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._31_  (.A(\u_usb_host.u_core.u_sie.u_crc5._00_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._01_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._02_ ));
 sky130_fd_sc_hd__xnor2_2 \u_usb_host.u_core.u_sie.u_crc5._32_  (.A(\u_usb_host.u_core.u_sie.token_q[11] ),
    .B(\u_usb_host.u_core.u_sie.token_q[8] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._03_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._33_  (.A(\u_usb_host.u_core.u_sie.token_q[10] ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._03_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._04_ ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc5._34_  (.A(net559),
    .B(net550),
    .X(\u_usb_host.u_core.u_sie.u_crc5._05_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._34__550  (.HI(net550));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._34__559  (.HI(net559));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._35_  (.A(\u_usb_host.u_core.u_sie.u_crc5._02_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._05_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._06_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._36_  (.A(\u_usb_host.u_core.u_sie.u_crc5._04_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._06_ ),
    .Y(\u_usb_host.u_core.u_sie.crc5_out_w[0] ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._37_  (.A(\u_usb_host.u_core.u_sie.token_q[12] ),
    .B(\u_usb_host.u_core.u_sie.token_q[6] ),
    .X(\u_usb_host.u_core.u_sie.u_crc5._07_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._38_  (.A(\u_usb_host.u_core.u_sie.token_q[11] ),
    .B(\u_usb_host.u_core.u_sie.token_q[9] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._08_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._39_  (.A(\u_usb_host.u_core.u_sie.u_crc5._07_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._08_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._09_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._40_  (.A(\u_usb_host.u_core.u_sie.token_q[15] ),
    .B(net551),
    .X(\u_usb_host.u_core.u_sie.u_crc5._10_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._40__551  (.HI(net551));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._41_  (.A(\u_usb_host.u_core.u_sie.u_crc5._05_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._10_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._11_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._42_  (.A(\u_usb_host.u_core.u_sie.u_crc5._09_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._11_ ),
    .Y(\u_usb_host.u_core.u_sie.crc5_out_w[1] ));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc5._43_  (.A(\u_usb_host.u_core.u_sie.token_q[13] ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._00_ ),
    .X(\u_usb_host.u_core.u_sie.u_crc5._12_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._44_  (.A(net554),
    .B(\u_usb_host.u_core.u_sie.u_crc5._12_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._13_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._44__554  (.HI(net554));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._45_  (.A(net552),
    .B(\u_usb_host.u_core.u_sie.u_crc5._03_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._14_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._45__552  (.HI(net552));
 sky130_fd_sc_hd__xor2_2 \u_usb_host.u_core.u_sie.u_crc5._46_  (.A(net557),
    .B(\u_usb_host.u_core.u_sie.token_q[7] ),
    .X(\u_usb_host.u_core.u_sie.u_crc5._15_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._46__557  (.HI(net557));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._47_  (.A(\u_usb_host.u_core.u_sie.token_q[5] ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._15_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._16_ ));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._48_  (.A(\u_usb_host.u_core.u_sie.token_q[12] ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._05_ ),
    .X(\u_usb_host.u_core.u_sie.u_crc5._17_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._49_  (.A(\u_usb_host.u_core.u_sie.u_crc5._16_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._17_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._18_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._50_  (.A(\u_usb_host.u_core.u_sie.u_crc5._14_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._18_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._19_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._51_  (.A(\u_usb_host.u_core.u_sie.u_crc5._13_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._19_ ),
    .Y(\u_usb_host.u_core.u_sie.crc5_out_w[2] ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._52_  (.A(net560),
    .B(\u_usb_host.u_core.u_sie.u_crc5._07_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._20_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._52__560  (.HI(net560));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._53_  (.A(\u_usb_host.u_core.u_sie.token_q[8] ),
    .B(net558),
    .X(\u_usb_host.u_core.u_sie.u_crc5._21_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._53__558  (.HI(net558));
 sky130_fd_sc_hd__xor2_1 \u_usb_host.u_core.u_sie.u_crc5._54_  (.A(\u_usb_host.u_core.u_sie.token_q[9] ),
    .B(net553),
    .X(\u_usb_host.u_core.u_sie.u_crc5._22_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._54__553  (.HI(net553));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._55_  (.A(\u_usb_host.u_core.u_sie.u_crc5._21_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._22_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._23_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._56_  (.A(\u_usb_host.u_core.u_sie.u_crc5._20_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._23_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._24_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._57_  (.A(\u_usb_host.u_core.u_sie.u_crc5._13_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._24_ ),
    .Y(\u_usb_host.u_core.u_sie.crc5_out_w[3] ));
 sky130_fd_sc_hd__xnor2_2 \u_usb_host.u_core.u_sie.u_crc5._58_  (.A(net561),
    .B(net555),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._25_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._58__555  (.HI(net555));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_core.u_sie.u_crc5._58__561  (.HI(net561));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._59_  (.A(\u_usb_host.u_core.u_sie.token_q[10] ),
    .B(\u_usb_host.u_core.u_sie.token_q[9] ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._26_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._60_  (.A(\u_usb_host.u_core.u_sie.u_crc5._25_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._26_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._27_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._61_  (.A(\u_usb_host.u_core.u_sie.u_crc5._12_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._27_ ),
    .Y(\u_usb_host.u_core.u_sie.u_crc5._28_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_core.u_sie.u_crc5._62_  (.A(\u_usb_host.u_core.u_sie.u_crc5._15_ ),
    .B(\u_usb_host.u_core.u_sie.u_crc5._28_ ),
    .Y(\u_usb_host.u_core.u_sie.crc5_out_w[4] ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._184_  (.A(net419),
    .Y(\u_usb_host.u_phy._051_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._185_  (.A(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .Y(\u_usb_host.u_phy._052_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._186_  (.A(\u_usb_host.u_phy.ones_count_q[0] ),
    .Y(\u_usb_host.u_phy._053_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._187_  (.A(\u_usb_host.u_core.u_sie.utmi_txvalid_o ),
    .Y(\u_usb_host.u_phy._054_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._188_  (.A(\u_usb_host.u_phy.send_eop_q ),
    .Y(\u_usb_host.u_phy._055_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._189_  (.A(\u_usb_host.u_phy.adjust_delayed_q ),
    .Y(\u_usb_host.u_phy._037_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_phy._190_  (.A(\u_usb_host.u_phy.usb_tx_dp_o ),
    .Y(\u_usb_host.u_phy._056_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._191__1  (.A(clknet_leaf_14_usb_clk),
    .Y(net564));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._192_  (.A(net418),
    .B(net417),
    .X(\u_usb_host.u_phy._057_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._193_  (.A(net421),
    .B(\u_usb_host.u_phy._057_ ),
    .Y(\u_usb_host.u_phy._046_ ));
 sky130_fd_sc_hd__nor4_2 \u_usb_host.u_phy._194_  (.A(net418),
    .B(net417),
    .C(\u_usb_host.u_phy.state_q[0] ),
    .D(net419),
    .Y(\u_usb_host.u_phy._058_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._195_  (.A(net117),
    .Y(\u_usb_host.u_phy._031_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._196_  (.A_N(\u_usb_host.u_phy.state_q[3] ),
    .B(net418),
    .X(\u_usb_host.u_phy._059_ ));
 sky130_fd_sc_hd__or3b_4 \u_usb_host.u_phy._197_  (.A(net421),
    .B(net419),
    .C_N(\u_usb_host.u_phy._059_ ),
    .X(\u_usb_host.u_phy._060_ ));
 sky130_fd_sc_hd__clkinv_2 \u_usb_host.u_phy._198_  (.A(\u_usb_host.u_phy._060_ ),
    .Y(\u_usb_host.u_core.u_sie.utmi_rxactive_i ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._199_  (.A(\u_usb_host.u_phy._053_ ),
    .B(\u_usb_host.u_phy.ones_count_q[1] ),
    .X(\u_usb_host.u_phy._061_ ));
 sky130_fd_sc_hd__nand3b_1 \u_usb_host.u_phy._200_  (.A_N(\u_usb_host.u_phy.ones_count_q[0] ),
    .B(\u_usb_host.u_phy.ones_count_q[1] ),
    .C(\u_usb_host.u_phy.ones_count_q[2] ),
    .Y(\u_usb_host.u_phy._062_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._201_  (.A(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .X(\u_usb_host.u_phy._063_ ));
 sky130_fd_sc_hd__nor3_2 \u_usb_host.u_phy._202_  (.A(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .C(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .Y(\u_usb_host.u_phy._064_ ));
 sky130_fd_sc_hd__or3_2 \u_usb_host.u_phy._203_  (.A(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .C(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .X(\u_usb_host.u_phy._065_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._204_  (.A_N(net418),
    .B(net417),
    .X(\u_usb_host.u_phy._066_ ));
 sky130_fd_sc_hd__nand2b_1 \u_usb_host.u_phy._205_  (.A_N(net418),
    .B(net417),
    .Y(\u_usb_host.u_phy._067_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._206_  (.A(net115),
    .B(\u_usb_host.u_phy._067_ ),
    .Y(\u_usb_host.u_phy._068_ ));
 sky130_fd_sc_hd__or4b_2 \u_usb_host.u_phy._207_  (.A(net418),
    .B(\u_usb_host.u_phy.state_q[0] ),
    .C(net420),
    .D_N(net417),
    .X(\u_usb_host.u_phy._069_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._208_  (.A(net115),
    .B(\u_usb_host.u_phy._069_ ),
    .Y(\u_usb_host.u_phy._070_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._209_  (.A(\u_usb_host.u_phy._062_ ),
    .B(\u_usb_host.u_phy._070_ ),
    .X(\u_usb_host.u_phy._071_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._210_  (.A(net421),
    .B(net419),
    .C(\u_usb_host.u_phy._059_ ),
    .X(\u_usb_host.u_phy._072_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._211_  (.A(net116),
    .B(\u_usb_host.u_phy._072_ ),
    .X(\u_usb_host.u_phy._073_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._212_  (.A(\u_usb_host.u_phy._060_ ),
    .B(\u_usb_host.u_phy._065_ ),
    .Y(\u_usb_host.u_phy._074_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._213_  (.A(\u_usb_host.u_core.u_sie.utmi_rxactive_i ),
    .B(\u_usb_host.u_phy._062_ ),
    .C(\u_usb_host.u_phy._064_ ),
    .X(\u_usb_host.u_phy._075_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._214_  (.A(net117),
    .B(\u_usb_host.u_phy._071_ ),
    .C(\u_usb_host.u_phy._073_ ),
    .D(\u_usb_host.u_phy._075_ ),
    .X(\u_usb_host.u_phy._047_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._215_  (.A(net421),
    .B(\u_usb_host.u_phy._051_ ),
    .Y(\u_usb_host.u_phy._076_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._216_  (.A_N(net419),
    .B(net421),
    .X(\u_usb_host.u_phy._077_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_phy._217_  (.A(net421),
    .B(net419),
    .Y(\u_usb_host.u_phy._078_ ));
 sky130_fd_sc_hd__or4bb_1 \u_usb_host.u_phy._218_  (.A(net418),
    .B(net417),
    .C_N(net421),
    .D_N(net420),
    .X(\u_usb_host.u_phy._079_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._219_  (.A(\u_usb_host.u_phy._079_ ),
    .Y(\u_usb_host.u_phy._080_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._220_  (.A(\u_usb_host.u_phy._058_ ),
    .B(\u_usb_host.u_phy._080_ ),
    .Y(\u_usb_host.u_phy._081_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._221_  (.A(net420),
    .B(\u_usb_host.u_phy._046_ ),
    .C(net116),
    .X(\u_usb_host.u_phy._082_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_phy._222_  (.A(\u_usb_host.u_phy._082_ ),
    .B(\u_usb_host.u_phy._047_ ),
    .C_N(\u_usb_host.u_phy._081_ ),
    .X(\u_usb_host.u_phy._043_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._223_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .Y(\u_usb_host.u_phy._083_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._224_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .X(\u_usb_host.u_phy._084_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._225_  (.A(\u_usb_host.u_phy.rxd_q ),
    .B(\u_usb_host.u_phy._084_ ),
    .X(\u_usb_host.u_phy.in_j_w ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_phy._226_  (.A(\u_usb_host.u_core.utmi_xcvrselect_o[1] ),
    .B(\u_usb_host.u_core.utmi_xcvrselect_o[0] ),
    .C(\u_usb_host.u_core.utmi_termselect_o ),
    .D(\u_usb_host.u_core.utmi_op_mode_o[0] ),
    .Y(\u_usb_host.u_phy._085_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_phy._227_  (.A1(\u_usb_host.u_core.utmi_op_mode_o[1] ),
    .A2(\u_usb_host.u_core.utmi_dppulldown_o ),
    .A3(\u_usb_host.u_core.utmi_dmpulldown_o ),
    .A4(\u_usb_host.u_phy._085_ ),
    .B1(net544),
    .X(\u_usb_host.u_phy._086_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_phy._227__544  (.LO(net544));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._228_  (.A(net418),
    .B(net417),
    .C(\u_usb_host.u_phy._077_ ),
    .D(\u_usb_host.u_phy._086_ ),
    .X(\u_usb_host.u_phy._087_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._229_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[2] ),
    .C(\u_usb_host.u_phy._065_ ),
    .D_N(\u_usb_host.u_phy.bit_count_q[0] ),
    .X(\u_usb_host.u_phy._088_ ));
 sky130_fd_sc_hd__o21ba_1 \u_usb_host.u_phy._230_  (.A1(\u_usb_host.u_phy.rx_dn_q ),
    .A2(\u_usb_host.u_phy.rx_dp_q ),
    .B1_N(\u_usb_host.u_phy.rxd_q ),
    .X(\u_usb_host.u_phy._089_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._231_  (.A(\u_usb_host.u_phy._064_ ),
    .B(\u_usb_host.u_phy._084_ ),
    .Y(\u_usb_host.u_phy._090_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._232_  (.A(net116),
    .B(\u_usb_host.u_phy._089_ ),
    .Y(\u_usb_host.u_phy._091_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_phy._233_  (.A1(net420),
    .A2(\u_usb_host.u_phy._046_ ),
    .A3(\u_usb_host.u_phy._088_ ),
    .A4(\u_usb_host.u_phy._091_ ),
    .B1(\u_usb_host.u_phy._087_ ),
    .X(\u_usb_host.u_phy._092_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._234_  (.A(\u_usb_host.u_phy.rx_dn_q ),
    .B(\u_usb_host.u_phy.rx_dp_q ),
    .C(net116),
    .X(\u_usb_host.u_phy._093_ ));
 sky130_fd_sc_hd__a211oi_1 \u_usb_host.u_phy._235_  (.A1(\u_usb_host.u_phy._064_ ),
    .A2(\u_usb_host.u_phy._083_ ),
    .B1(\u_usb_host.u_phy._093_ ),
    .C1(\u_usb_host.u_phy._060_ ),
    .Y(\u_usb_host.u_phy._094_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._236_  (.A(\u_usb_host.u_phy.state_q[0] ),
    .B(net420),
    .C(\u_usb_host.u_phy._066_ ),
    .X(\u_usb_host.u_phy._095_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._237_  (.A(\u_usb_host.u_core.u_sie.utmi_txvalid_o ),
    .B(\u_usb_host.u_phy._086_ ),
    .X(\u_usb_host.u_phy._096_ ));
 sky130_fd_sc_hd__nor3_1 \u_usb_host.u_phy._238_  (.A(\u_usb_host.u_phy._031_ ),
    .B(\u_usb_host.u_phy._089_ ),
    .C(\u_usb_host.u_phy._096_ ),
    .Y(\u_usb_host.u_phy._097_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._239_  (.A(\u_usb_host.u_phy._067_ ),
    .B(\u_usb_host.u_phy._078_ ),
    .Y(\u_usb_host.u_phy._098_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._240_  (.A(net418),
    .B(net417),
    .C(net419),
    .X(\u_usb_host.u_phy._099_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._241_  (.A1(\u_usb_host.u_phy._054_ ),
    .A2(\u_usb_host.u_phy.send_eop_q ),
    .B1(\u_usb_host.u_phy._062_ ),
    .X(\u_usb_host.u_phy._100_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._242_  (.A(\u_usb_host.u_phy._069_ ),
    .B(\u_usb_host.u_phy._100_ ),
    .Y(\u_usb_host.u_phy._101_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._243_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .Y(\u_usb_host.u_phy._102_ ));
 sky130_fd_sc_hd__nand3_2 \u_usb_host.u_phy._244_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .C(\u_usb_host.u_phy.bit_count_q[2] ),
    .Y(\u_usb_host.u_phy._103_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._245_  (.A(\u_usb_host.u_phy._080_ ),
    .B(\u_usb_host.u_phy._090_ ),
    .X(\u_usb_host.u_phy._104_ ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_phy._246_  (.A1(net115),
    .A2(\u_usb_host.u_phy._095_ ),
    .B1(\u_usb_host.u_phy._099_ ),
    .C1(\u_usb_host.u_phy._104_ ),
    .D1(\u_usb_host.u_phy._094_ ),
    .X(\u_usb_host.u_phy._105_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_phy._247_  (.A1(\u_usb_host.u_phy._065_ ),
    .A2(\u_usb_host.u_phy._098_ ),
    .B1_N(\u_usb_host.u_phy._069_ ),
    .X(\u_usb_host.u_phy._106_ ));
 sky130_fd_sc_hd__o32a_1 \u_usb_host.u_phy._248_  (.A1(\u_usb_host.u_phy._065_ ),
    .A2(\u_usb_host.u_phy._101_ ),
    .A3(\u_usb_host.u_phy._103_ ),
    .B1(\u_usb_host.u_phy._106_ ),
    .B2(\u_usb_host.u_phy._072_ ),
    .X(\u_usb_host.u_phy._107_ ));
 sky130_fd_sc_hd__nor4_1 \u_usb_host.u_phy._249_  (.A(\u_usb_host.u_phy._092_ ),
    .B(\u_usb_host.u_phy._097_ ),
    .C(\u_usb_host.u_phy._105_ ),
    .D(\u_usb_host.u_phy._107_ ),
    .Y(\u_usb_host.u_phy._042_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._250_  (.A(\u_usb_host.u_core.u_sie.utmi_txvalid_o ),
    .B(\u_usb_host.u_phy._069_ ),
    .Y(\u_usb_host.u_phy._030_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._251_  (.A1(\u_usb_host.u_phy._066_ ),
    .A2(\u_usb_host.u_phy._076_ ),
    .B1(\u_usb_host.u_phy._030_ ),
    .X(\u_usb_host.u_phy._045_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._252_  (.A(net685),
    .B(\u_usb_host.u_phy.rxd0_q ),
    .X(\u_usb_host.u_phy._022_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._253_  (.A(\u_usb_host.u_phy.rxd1_q ),
    .B(\u_usb_host.u_phy.rxd0_q ),
    .Y(\u_usb_host.u_phy._108_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._254_  (.A(\u_usb_host.u_phy._022_ ),
    .B(\u_usb_host.u_phy._108_ ),
    .X(\u_usb_host.u_phy._041_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_phy._255_  (.A(net117),
    .B(\u_usb_host.u_phy._070_ ),
    .C(\u_usb_host.u_phy._074_ ),
    .X(\u_usb_host.u_phy._040_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._256_  (.A(\u_usb_host.u_phy.rx_dn1_q ),
    .B(\u_usb_host.u_phy.rx_dn0_q ),
    .X(\u_usb_host.u_phy._017_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._257_  (.A(\u_usb_host.u_phy.rx_dn1_q ),
    .B(\u_usb_host.u_phy.rx_dn0_q ),
    .Y(\u_usb_host.u_phy._109_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._258_  (.A(\u_usb_host.u_phy._017_ ),
    .B(\u_usb_host.u_phy._109_ ),
    .X(\u_usb_host.u_phy._039_ ));
 sky130_fd_sc_hd__and2_1 \u_usb_host.u_phy._259_  (.A(net686),
    .B(\u_usb_host.u_phy.rx_dp0_q ),
    .X(\u_usb_host.u_phy._018_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._260_  (.A(\u_usb_host.u_phy.rx_dp1_q ),
    .B(\u_usb_host.u_phy.rx_dp0_q ),
    .Y(\u_usb_host.u_phy._110_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._261_  (.A(\u_usb_host.u_phy._018_ ),
    .B(\u_usb_host.u_phy._110_ ),
    .X(\u_usb_host.u_phy._038_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._266_  (.A(net117),
    .B(net116),
    .X(\u_usb_host.u_phy._036_ ));
 sky130_fd_sc_hd__or4bb_1 \u_usb_host.u_phy._267_  (.A(net421),
    .B(net419),
    .C_N(net418),
    .D_N(net417),
    .X(\u_usb_host.u_phy._113_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._268_  (.A1(net115),
    .A2(\u_usb_host.u_phy._113_ ),
    .B1(\u_usb_host.u_phy._031_ ),
    .Y(\u_usb_host.u_phy._034_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._269_  (.A(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .B(\u_usb_host.u_phy._062_ ),
    .Y(\u_usb_host.u_phy._114_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._270_  (.A(\u_usb_host.u_phy._114_ ),
    .Y(\u_usb_host.u_phy._115_ ));
 sky130_fd_sc_hd__a311o_1 \u_usb_host.u_phy._271_  (.A1(\u_usb_host.u_phy.state_q[2] ),
    .A2(\u_usb_host.u_phy.state_q[3] ),
    .A3(\u_usb_host.u_phy._077_ ),
    .B1(\u_usb_host.u_phy._034_ ),
    .C1(\u_usb_host.u_phy._068_ ),
    .X(\u_usb_host.u_phy._116_ ));
 sky130_fd_sc_hd__o32a_1 \u_usb_host.u_phy._272_  (.A1(net419),
    .A2(\u_usb_host.u_phy._067_ ),
    .A3(\u_usb_host.u_phy._114_ ),
    .B1(\u_usb_host.u_phy._116_ ),
    .B2(\u_usb_host.u_phy._073_ ),
    .X(\u_usb_host.u_phy._033_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._273_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .C(\u_usb_host.u_phy.bit_count_q[2] ),
    .D(\u_usb_host.u_phy._075_ ),
    .X(\u_usb_host.u_phy._021_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._274_  (.A(net419),
    .B(\u_usb_host.u_phy.usb_tx_dn_o ),
    .C(net115),
    .D(\u_usb_host.u_phy._067_ ),
    .X(\u_usb_host.u_phy._117_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._275_  (.A0(\u_usb_host.u_phy._117_ ),
    .A1(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .S(\u_usb_host.u_phy._073_ ),
    .X(\u_usb_host.u_phy._118_ ));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_phy._276_  (.A(\u_usb_host.u_phy._118_ ),
    .Y(\u_usb_host.u_phy._015_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._277_  (.A(\u_usb_host.u_phy._075_ ),
    .B(\u_usb_host.u_phy._103_ ),
    .Y(\u_usb_host.u_phy._119_ ));
 sky130_fd_sc_hd__or2_2 \u_usb_host.u_phy._278_  (.A(\u_usb_host.u_phy._075_ ),
    .B(\u_usb_host.u_phy._103_ ),
    .X(\u_usb_host.u_phy._120_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._279_  (.A(\u_usb_host.u_core.u_sie.utmi_data_i[1] ),
    .B(\u_usb_host.u_phy._119_ ),
    .X(\u_usb_host.u_phy._121_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._280_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_o[0] ),
    .A2(\u_usb_host.u_phy._120_ ),
    .B1(\u_usb_host.u_phy._121_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._004_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._281_  (.A0(\u_usb_host.u_core.u_sie.utmi_data_o[1] ),
    .A1(\u_usb_host.u_core.u_sie.utmi_data_i[2] ),
    .S(\u_usb_host.u_phy._120_ ),
    .X(\u_usb_host.u_phy._122_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._282_  (.A(net117),
    .B(\u_usb_host.u_phy._122_ ),
    .X(\u_usb_host.u_phy._005_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._283_  (.A(\u_usb_host.u_core.u_sie.utmi_data_i[3] ),
    .B(\u_usb_host.u_phy._119_ ),
    .X(\u_usb_host.u_phy._123_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._284_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_o[2] ),
    .A2(\u_usb_host.u_phy._120_ ),
    .B1(\u_usb_host.u_phy._123_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._006_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._285_  (.A0(\u_usb_host.u_core.u_sie.utmi_data_o[3] ),
    .A1(\u_usb_host.u_core.u_sie.utmi_data_i[4] ),
    .S(\u_usb_host.u_phy._120_ ),
    .X(\u_usb_host.u_phy._124_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._286_  (.A(net117),
    .B(\u_usb_host.u_phy._124_ ),
    .X(\u_usb_host.u_phy._007_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._287_  (.A(\u_usb_host.u_core.u_sie.utmi_data_i[5] ),
    .B(\u_usb_host.u_phy._119_ ),
    .X(\u_usb_host.u_phy._125_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._288_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_o[4] ),
    .A2(\u_usb_host.u_phy._120_ ),
    .B1(\u_usb_host.u_phy._125_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._008_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._289_  (.A0(\u_usb_host.u_core.u_sie.utmi_data_o[5] ),
    .A1(\u_usb_host.u_core.u_sie.utmi_data_i[6] ),
    .S(\u_usb_host.u_phy._120_ ),
    .X(\u_usb_host.u_phy._126_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._290_  (.A(net117),
    .B(\u_usb_host.u_phy._126_ ),
    .X(\u_usb_host.u_phy._009_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._291_  (.A(\u_usb_host.u_core.u_sie.utmi_data_i[7] ),
    .B(\u_usb_host.u_phy._119_ ),
    .X(\u_usb_host.u_phy._127_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._292_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_o[6] ),
    .A2(\u_usb_host.u_phy._120_ ),
    .B1(\u_usb_host.u_phy._127_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._010_ ));
 sky130_fd_sc_hd__a31o_1 \u_usb_host.u_phy._293_  (.A1(\u_usb_host.u_phy.rxd_q ),
    .A2(\u_usb_host.u_phy.rxd_last_j_q ),
    .A3(\u_usb_host.u_phy._084_ ),
    .B1(net115),
    .X(\u_usb_host.u_phy._128_ ));
 sky130_fd_sc_hd__o21bai_4 \u_usb_host.u_phy._294_  (.A1(net671),
    .A2(\u_usb_host.u_phy.in_j_w ),
    .B1_N(\u_usb_host.u_phy._128_ ),
    .Y(\u_usb_host.u_phy._129_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._295_  (.A(\u_usb_host.u_phy._119_ ),
    .B(\u_usb_host.u_phy._129_ ),
    .X(\u_usb_host.u_phy._130_ ));
 sky130_fd_sc_hd__o211a_1 \u_usb_host.u_phy._296_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_o[7] ),
    .A2(\u_usb_host.u_phy._120_ ),
    .B1(\u_usb_host.u_phy._130_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._011_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._297_  (.A_N(\u_usb_host.u_phy.bit_count_q[0] ),
    .B(\u_usb_host.u_phy._081_ ),
    .X(\u_usb_host.u_phy._001_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._298_  (.A(\u_usb_host.u_phy.bit_count_q[1] ),
    .B(\u_usb_host.u_phy.bit_count_q[0] ),
    .X(\u_usb_host.u_phy._131_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._299_  (.A(\u_usb_host.u_phy._081_ ),
    .B(\u_usb_host.u_phy._102_ ),
    .C(\u_usb_host.u_phy._131_ ),
    .X(\u_usb_host.u_phy._002_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._300_  (.A1(\u_usb_host.u_phy.bit_count_q[1] ),
    .A2(\u_usb_host.u_phy.bit_count_q[0] ),
    .B1(\u_usb_host.u_phy.bit_count_q[2] ),
    .X(\u_usb_host.u_phy._132_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._301_  (.A(\u_usb_host.u_phy._081_ ),
    .B(\u_usb_host.u_phy._103_ ),
    .C(\u_usb_host.u_phy._132_ ),
    .X(\u_usb_host.u_phy._003_ ));
 sky130_fd_sc_hd__o221a_1 \u_usb_host.u_phy._302_  (.A1(\u_usb_host.u_phy._074_ ),
    .A2(\u_usb_host.u_phy._115_ ),
    .B1(\u_usb_host.u_phy._129_ ),
    .B2(\u_usb_host.u_phy._060_ ),
    .C1(\u_usb_host.u_phy._053_ ),
    .X(\u_usb_host.u_phy._133_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._303_  (.A(net117),
    .B(\u_usb_host.u_phy._133_ ),
    .X(\u_usb_host.u_phy._012_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._304_  (.A_N(\u_usb_host.u_phy.ones_count_q[1] ),
    .B(\u_usb_host.u_phy.ones_count_q[0] ),
    .X(\u_usb_host.u_phy._134_ ));
 sky130_fd_sc_hd__o221a_1 \u_usb_host.u_phy._305_  (.A1(\u_usb_host.u_phy._074_ ),
    .A2(\u_usb_host.u_phy._115_ ),
    .B1(\u_usb_host.u_phy._129_ ),
    .B2(\u_usb_host.u_phy._060_ ),
    .C1(\u_usb_host.u_phy._031_ ),
    .X(\u_usb_host.u_phy._135_ ));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_phy._306_  (.A1(\u_usb_host.u_phy._061_ ),
    .A2(\u_usb_host.u_phy._134_ ),
    .B1(\u_usb_host.u_phy._135_ ),
    .X(\u_usb_host.u_phy._013_ ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._307_  (.A1(\u_usb_host.u_phy.ones_count_q[0] ),
    .A2(\u_usb_host.u_phy.ones_count_q[1] ),
    .B1(\u_usb_host.u_phy.ones_count_q[2] ),
    .X(\u_usb_host.u_phy._136_ ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_phy._308_  (.A(\u_usb_host.u_phy.ones_count_q[2] ),
    .B(\u_usb_host.u_phy.ones_count_q[0] ),
    .C(\u_usb_host.u_phy.ones_count_q[1] ),
    .Y(\u_usb_host.u_phy._137_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._309_  (.A(\u_usb_host.u_phy._135_ ),
    .B(\u_usb_host.u_phy._136_ ),
    .C(\u_usb_host.u_phy._137_ ),
    .X(\u_usb_host.u_phy._014_ ));
 sky130_fd_sc_hd__xnor2_1 \u_usb_host.u_phy._310_  (.A(net580),
    .B(\u_usb_host.u_phy.in_j_w ),
    .Y(\u_usb_host.u_phy._138_ ));
 sky130_fd_sc_hd__nor3_2 \u_usb_host.u_phy._311_  (.A(\u_usb_host.u_phy.state_q[3] ),
    .B(\u_usb_host.u_phy._072_ ),
    .C(\u_usb_host.u_phy._138_ ),
    .Y(\u_usb_host.u_phy._139_ ));
 sky130_fd_sc_hd__o31ai_1 \u_usb_host.u_phy._312_  (.A1(\u_usb_host.u_phy._052_ ),
    .A2(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .A3(\u_usb_host.u_phy._139_ ),
    .B1(net115),
    .Y(\u_usb_host.u_phy._048_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._313_  (.A(\u_usb_host.u_phy.sample_cnt_q[1] ),
    .B(\u_usb_host.u_phy.sample_cnt_q[0] ),
    .Y(\u_usb_host.u_phy._140_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._314_  (.A(\u_usb_host.u_phy._063_ ),
    .B(\u_usb_host.u_phy._140_ ),
    .Y(\u_usb_host.u_phy._141_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._315_  (.A(\u_usb_host.u_phy._139_ ),
    .B(\u_usb_host.u_phy._141_ ),
    .Y(\u_usb_host.u_phy._049_ ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_phy._316_  (.A0(\u_usb_host.u_phy._140_ ),
    .A1(\u_usb_host.u_phy._141_ ),
    .S(\u_usb_host.u_phy.sample_cnt_q[2] ),
    .X(\u_usb_host.u_phy._142_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._317_  (.A(\u_usb_host.u_phy._139_ ),
    .B(\u_usb_host.u_phy._142_ ),
    .Y(\u_usb_host.u_phy._050_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._318_  (.A(\u_usb_host.u_phy._037_ ),
    .B(net116),
    .C(\u_usb_host.u_phy._139_ ),
    .X(\u_usb_host.u_phy._000_ ));
 sky130_fd_sc_hd__nand2_1 \u_usb_host.u_phy._333_  (.A(net117),
    .B(\u_usb_host.u_phy._096_ ),
    .Y(\u_usb_host.u_phy._019_ ));
 sky130_fd_sc_hd__mux2_2 \u_usb_host.u_phy._334_  (.A0(\u_usb_host.u_phy.usb_tx_dp_o ),
    .A1(\u_usb_host.u_phy.rx_dp_q ),
    .S(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(\u_usb_host.u_core.u_sie.utmi_linestate_i[0] ));
 sky130_fd_sc_hd__mux2_2 \u_usb_host.u_phy._335_  (.A0(\u_usb_host.u_phy.usb_tx_dn_o ),
    .A1(\u_usb_host.u_phy.rx_dn_q ),
    .S(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(\u_usb_host.u_core.u_sie.utmi_linestate_i[1] ));
 sky130_fd_sc_hd__nand3_1 \u_usb_host.u_phy._336_  (.A(\u_usb_host.u_phy.ones_count_q[2] ),
    .B(\u_usb_host.u_phy._129_ ),
    .C(\u_usb_host.u_phy._134_ ),
    .Y(\u_usb_host.u_phy._150_ ));
 sky130_fd_sc_hd__or3b_1 \u_usb_host.u_phy._337_  (.A(net417),
    .B(net116),
    .C_N(\u_usb_host.u_phy._077_ ),
    .X(\u_usb_host.u_phy._151_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._338_  (.A(net117),
    .B(\u_usb_host.u_phy._099_ ),
    .Y(\u_usb_host.u_phy._152_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_phy._339_  (.A1(net421),
    .A2(\u_usb_host.u_phy._051_ ),
    .A3(\u_usb_host.u_phy._067_ ),
    .B1(\u_usb_host.u_phy._151_ ),
    .C1(\u_usb_host.u_phy._152_ ),
    .X(\u_usb_host.u_phy._153_ ));
 sky130_fd_sc_hd__or4b_1 \u_usb_host.u_phy._340_  (.A(\u_usb_host.u_phy._057_ ),
    .B(net115),
    .C(\u_usb_host.u_phy._078_ ),
    .D_N(\u_usb_host.u_phy._089_ ),
    .X(\u_usb_host.u_phy._154_ ));
 sky130_fd_sc_hd__o311a_1 \u_usb_host.u_phy._341_  (.A1(\u_usb_host.u_phy._060_ ),
    .A2(net115),
    .A3(\u_usb_host.u_phy._084_ ),
    .B1(\u_usb_host.u_phy._153_ ),
    .C1(\u_usb_host.u_phy._154_ ),
    .X(\u_usb_host.u_phy._155_ ));
 sky130_fd_sc_hd__o21ai_1 \u_usb_host.u_phy._342_  (.A1(\u_usb_host.u_phy._069_ ),
    .A2(\u_usb_host.u_phy._150_ ),
    .B1(\u_usb_host.u_phy._155_ ),
    .Y(\u_usb_host.u_phy.next_state_r[0] ));
 sky130_fd_sc_hd__a31oi_1 \u_usb_host.u_phy._343_  (.A1(\u_usb_host.u_phy.ones_count_q[2] ),
    .A2(\u_usb_host.u_phy._129_ ),
    .A3(\u_usb_host.u_phy._134_ ),
    .B1(\u_usb_host.u_phy._069_ ),
    .Y(\u_usb_host.u_phy._156_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._344_  (.A(\u_usb_host.u_phy._059_ ),
    .B(net115),
    .C(\u_usb_host.u_phy._076_ ),
    .X(\u_usb_host.u_phy._157_ ));
 sky130_fd_sc_hd__and4_1 \u_usb_host.u_phy._345_  (.A(\u_usb_host.u_phy._059_ ),
    .B(net116),
    .C(\u_usb_host.u_phy._077_ ),
    .D(\u_usb_host.u_phy._083_ ),
    .X(\u_usb_host.u_phy._158_ ));
 sky130_fd_sc_hd__a21bo_1 \u_usb_host.u_phy._346_  (.A1(\u_usb_host.u_phy._080_ ),
    .A2(\u_usb_host.u_phy._091_ ),
    .B1_N(\u_usb_host.u_phy._154_ ),
    .X(\u_usb_host.u_phy._159_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._347_  (.A(\u_usb_host.u_phy._098_ ),
    .B(\u_usb_host.u_phy._157_ ),
    .C(\u_usb_host.u_phy._158_ ),
    .D(\u_usb_host.u_phy._159_ ),
    .X(\u_usb_host.u_phy._160_ ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._348_  (.A(\u_usb_host.u_phy._089_ ),
    .B(\u_usb_host.u_phy._152_ ),
    .Y(\u_usb_host.u_phy._161_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_phy._349_  (.A1(\u_usb_host.u_core.u_sie.utmi_txvalid_o ),
    .A2(\u_usb_host.u_phy._161_ ),
    .B1(\u_usb_host.u_phy._160_ ),
    .C1(\u_usb_host.u_phy._156_ ),
    .X(\u_usb_host.u_phy.next_state_r[1] ));
 sky130_fd_sc_hd__nor2_1 \u_usb_host.u_phy._350_  (.A(net116),
    .B(\u_usb_host.u_phy._113_ ),
    .Y(\u_usb_host.u_phy._162_ ));
 sky130_fd_sc_hd__o2111a_1 \u_usb_host.u_phy._351_  (.A1(net421),
    .A2(net116),
    .B1(\u_usb_host.u_phy._090_ ),
    .C1(\u_usb_host.u_phy._051_ ),
    .D1(\u_usb_host.u_phy._059_ ),
    .X(\u_usb_host.u_phy._163_ ));
 sky130_fd_sc_hd__or4_1 \u_usb_host.u_phy._352_  (.A(\u_usb_host.u_phy._095_ ),
    .B(\u_usb_host.u_phy._157_ ),
    .C(\u_usb_host.u_phy._162_ ),
    .D(\u_usb_host.u_phy._163_ ),
    .X(\u_usb_host.u_phy._164_ ));
 sky130_fd_sc_hd__a41o_1 \u_usb_host.u_phy._353_  (.A1(net595),
    .A2(\u_usb_host.u_phy._064_ ),
    .A3(\u_usb_host.u_phy._080_ ),
    .A4(\u_usb_host.u_phy._089_ ),
    .B1(\u_usb_host.u_phy._161_ ),
    .X(\u_usb_host.u_phy._165_ ));
 sky130_fd_sc_hd__or2_1 \u_usb_host.u_phy._354_  (.A(\u_usb_host.u_phy._164_ ),
    .B(\u_usb_host.u_phy._165_ ),
    .X(\u_usb_host.u_phy.next_state_r[2] ));
 sky130_fd_sc_hd__a2111o_1 \u_usb_host.u_phy._355_  (.A1(\u_usb_host.u_phy._054_ ),
    .A2(\u_usb_host.u_phy._161_ ),
    .B1(\u_usb_host.u_phy._162_ ),
    .C1(\u_usb_host.u_phy._066_ ),
    .D1(\u_usb_host.u_phy._072_ ),
    .X(\u_usb_host.u_phy.next_state_r[3] ));
 sky130_fd_sc_hd__a21o_1 \u_usb_host.u_phy._356_  (.A1(\u_usb_host.u_phy._055_ ),
    .A2(\u_usb_host.u_phy._071_ ),
    .B1(\u_usb_host.u_phy._073_ ),
    .X(\u_usb_host.u_phy._166_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_phy._357_  (.A_N(\u_usb_host.u_phy._103_ ),
    .B(\u_usb_host.u_phy._166_ ),
    .X(\u_usb_host.u_phy._032_ ));
 sky130_fd_sc_hd__or3_1 \u_usb_host.u_phy._358_  (.A(\u_usb_host.u_phy.sync_j_detected_q ),
    .B(\u_usb_host.u_phy._079_ ),
    .C(\u_usb_host.u_phy._091_ ),
    .X(\u_usb_host.u_phy._167_ ));
 sky130_fd_sc_hd__nand3b_1 \u_usb_host.u_phy._359_  (.A_N(\u_usb_host.u_phy._093_ ),
    .B(\u_usb_host.u_phy._137_ ),
    .C(\u_usb_host.u_phy._167_ ),
    .Y(\u_usb_host.u_phy._020_ ));
 sky130_fd_sc_hd__and3_1 \u_usb_host.u_phy._360_  (.A(\u_usb_host.u_phy._051_ ),
    .B(\u_usb_host.u_phy._056_ ),
    .C(\u_usb_host.u_phy._068_ ),
    .X(\u_usb_host.u_phy._168_ ));
 sky130_fd_sc_hd__a211o_1 \u_usb_host.u_phy._361_  (.A1(\u_usb_host.u_core.u_sie.utmi_data_i[0] ),
    .A2(\u_usb_host.u_phy._073_ ),
    .B1(\u_usb_host.u_phy._034_ ),
    .C1(\u_usb_host.u_phy._168_ ),
    .X(\u_usb_host.u_phy._016_ ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_phy._369_  (.CLK(\u_usb_host.u_phy._170_ ),
    .D(\u_usb_host.u_phy._019_ ),
    .SET_B(net391),
    .Q(\u_usb_host.u_phy.usb_tx_oen_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._370_  (.CLK(\u_usb_host.u_phy._172_ ),
    .D(\u_usb_host.u_phy.in_j_w ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_phy.rxd_last_j_q ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_phy._371_  (.CLK(\u_usb_host.u_phy._183_ ),
    .D(\u_usb_host.u_phy._016_ ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_phy.usb_tx_dp_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._372_  (.CLK(\u_usb_host.u_phy._181_ ),
    .D(\u_usb_host.u_phy._031_ ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.sync_j_detected_q ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_phy._373_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._004_ ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._374_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._005_ ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._375_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._006_ ),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._376_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._007_ ),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._377_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._008_ ),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[4] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._378_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._009_ ),
    .RESET_B(net407),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[5] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._379_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._010_ ),
    .RESET_B(net405),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[6] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._380_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._182_ ),
    .D(\u_usb_host.u_phy._011_ ),
    .RESET_B(net408),
    .Q(\u_usb_host.u_core.u_sie.utmi_data_i[7] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._381_  (.CLK(\u_usb_host.u_phy._174_ ),
    .D(\u_usb_host.u_phy._018_ ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dp_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._382_  (.CLK(\u_usb_host.u_phy._169_ ),
    .D(\u_usb_host.u_phy._015_ ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_phy.usb_tx_dn_o ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._383_  (.CLK(\u_usb_host.u_phy._175_ ),
    .D(\u_usb_host.u_phy._017_ ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dn_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._384_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._173_ ),
    .D(\u_usb_host.u_phy._048_ ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.sample_cnt_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._385_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._173_ ),
    .D(\u_usb_host.u_phy._049_ ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.sample_cnt_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._386_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._173_ ),
    .D(\u_usb_host.u_phy._050_ ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.sample_cnt_q[2] ));
 sky130_fd_sc_hd__dfstp_1 \u_usb_host.u_phy._387_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._176_ ),
    .D(\u_usb_host.u_phy._012_ ),
    .SET_B(net395),
    .Q(\u_usb_host.u_phy.ones_count_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._388_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._176_ ),
    .D(\u_usb_host.u_phy._013_ ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.ones_count_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._389_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._176_ ),
    .D(\u_usb_host.u_phy._014_ ),
    .RESET_B(net409),
    .Q(\u_usb_host.u_phy.ones_count_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._390_  (.CLK(\u_usb_host.u_phy._177_ ),
    .D(\u_usb_host.u_phy._022_ ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rxd_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._391_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy.next_state_r[0] ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.state_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._392_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy.next_state_r[1] ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.state_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._393_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy.next_state_r[2] ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.state_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._394_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._178_ ),
    .D(\u_usb_host.u_phy.next_state_r[3] ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.state_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._395_  (.CLK(\u_usb_host.u_phy._180_ ),
    .D(\u_usb_host.u_phy._030_ ),
    .RESET_B(net395),
    .Q(\u_usb_host.u_phy.send_eop_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._396_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._179_ ),
    .D(\u_usb_host.u_phy._001_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_phy.bit_count_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._397_  (.CLK(\clknet_1_0__leaf_u_usb_host.u_phy._179_ ),
    .D(\u_usb_host.u_phy._002_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_phy.bit_count_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._398_  (.CLK(\clknet_1_1__leaf_u_usb_host.u_phy._179_ ),
    .D(\u_usb_host.u_phy._003_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_phy.bit_count_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._399_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_dp_i ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.rx_dp_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._400_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_dn_i ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dn_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._401_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy.usb_rx_rcv_i ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.rxd_ms ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._402_  (.CLK(clknet_leaf_10_usb_clk),
    .D(net683),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dp0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._403_  (.CLK(clknet_leaf_9_usb_clk),
    .D(net647),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dn0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._404_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy.rx_dp0_q ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dp1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._405_  (.CLK(clknet_leaf_9_usb_clk),
    .D(\u_usb_host.u_phy.rx_dn0_q ),
    .RESET_B(net389),
    .Q(\u_usb_host.u_phy.rx_dn1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._406_  (.CLK(clknet_leaf_10_usb_clk),
    .D(net678),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.rxd0_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._407_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy.rxd0_q ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.rxd1_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._408_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_phy._020_ ),
    .RESET_B(net391),
    .Q(\u_usb_host.u_core.utmi_rxerror_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._409_  (.CLK(clknet_leaf_11_usb_clk),
    .D(\u_usb_host.u_phy.in_j_w ),
    .RESET_B(net392),
    .Q(\u_usb_host.u_phy.rxd_last_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._410_  (.CLK(clknet_leaf_10_usb_clk),
    .D(\u_usb_host.u_phy._000_ ),
    .RESET_B(net390),
    .Q(\u_usb_host.u_phy.adjust_delayed_q ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_phy._411_  (.CLK(clknet_leaf_15_usb_clk),
    .D(\u_usb_host.u_phy._021_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.utmi_rxvalid_i ));
 sky130_fd_sc_hd__dfrtp_2 \u_usb_host.u_phy._412_  (.CLK(clknet_leaf_14_usb_clk),
    .D(\u_usb_host.u_phy._032_ ),
    .RESET_B(net406),
    .Q(\u_usb_host.u_core.u_sie.utmi_txready_i ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._413_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_phy._033_ ),
    .GCLK(\u_usb_host.u_phy._169_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._414_  (.CLK(clknet_leaf_10_usb_clk),
    .GATE(\u_usb_host.u_phy._034_ ),
    .GCLK(\u_usb_host.u_phy._170_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._416_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_phy._036_ ),
    .GCLK(\u_usb_host.u_phy._172_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._417_  (.CLK(clknet_leaf_10_usb_clk),
    .GATE(\u_usb_host.u_phy._037_ ),
    .GCLK(\u_usb_host.u_phy._173_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._418_  (.CLK(clknet_leaf_10_usb_clk),
    .GATE(\u_usb_host.u_phy._038_ ),
    .GCLK(\u_usb_host.u_phy._174_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._419_  (.CLK(clknet_leaf_9_usb_clk),
    .GATE(\u_usb_host.u_phy._039_ ),
    .GCLK(\u_usb_host.u_phy._175_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._420_  (.CLK(clknet_leaf_14_usb_clk),
    .GATE(\u_usb_host.u_phy._040_ ),
    .GCLK(\u_usb_host.u_phy._176_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._421_  (.CLK(clknet_leaf_10_usb_clk),
    .GATE(\u_usb_host.u_phy._041_ ),
    .GCLK(\u_usb_host.u_phy._177_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._422_  (.CLK(clknet_leaf_12_usb_clk),
    .GATE(\u_usb_host.u_phy._042_ ),
    .GCLK(\u_usb_host.u_phy._178_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._423_  (.CLK(clknet_leaf_14_usb_clk),
    .GATE(\u_usb_host.u_phy._043_ ),
    .GCLK(\u_usb_host.u_phy._179_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._424_  (.CLK(net564),
    .GATE(\u_usb_host.u_phy._045_ ),
    .GCLK(\u_usb_host.u_phy._180_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._425_  (.CLK(clknet_leaf_14_usb_clk),
    .GATE(\u_usb_host.u_phy._046_ ),
    .GCLK(\u_usb_host.u_phy._181_ ));
 sky130_fd_sc_hd__dlclkp_2 \u_usb_host.u_phy._426_  (.CLK(clknet_leaf_15_usb_clk),
    .GATE(\u_usb_host.u_phy._047_ ),
    .GCLK(\u_usb_host.u_phy._182_ ));
 sky130_fd_sc_hd__dlclkp_1 \u_usb_host.u_phy._427_  (.CLK(clknet_leaf_11_usb_clk),
    .GATE(\u_usb_host.u_phy._033_ ),
    .GCLK(\u_usb_host.u_phy._183_ ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_usb_rst._1_  (.CLK(clknet_leaf_0_usb_clk),
    .D(net562),
    .RESET_B(net46),
    .Q(\u_usb_host.u_usb_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_rst._1__562  (.HI(net562));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_usb_rst._2_  (.CLK(clknet_leaf_0_usb_clk),
    .D(net648),
    .RESET_B(net46),
    .Q(\u_usb_host.u_usb_rst.in_data_2s ));
 sky130_fd_sc_hd__mux2_4 \u_usb_host.u_usb_rst.u_buf.genblk1.u_mux  (.A0(net573),
    .A1(net46),
    .S(net545),
    .X(\u_usb_host.u_async_wb.u_cmd_if.rd_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_rst.u_buf.genblk1.u_mux_545  (.LO(net545));
 sky130_fd_sc_hd__inv_2 \u_usb_host.u_usb_xcvr._2_  (.A(\u_usb_host.u_phy.usb_tx_dn_o ),
    .Y(\u_usb_host.u_usb_xcvr._1_ ));
 sky130_fd_sc_hd__and2b_1 \u_usb_host.u_usb_xcvr._3_  (.A_N(net44),
    .B(net45),
    .X(\u_usb_host.u_phy.usb_rx_rcv_i ));
 sky130_fd_sc_hd__nor2_2 \u_usb_host.u_usb_xcvr._4_  (.A(\u_usb_host.u_phy.usb_tx_dp_o ),
    .B(net547),
    .Y(\u_usb_host.u_usb_xcvr._0_ ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._4__547  (.HI(net547));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_usb_xcvr._5_  (.A0(net548),
    .A1(\u_usb_host.u_usb_xcvr._0_ ),
    .S(\u_usb_host.u_usb_xcvr._1_ ),
    .X(net82));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._5__548  (.HI(net548));
 sky130_fd_sc_hd__o21a_1 \u_usb_host.u_usb_xcvr._6_  (.A1(\u_usb_host.u_usb_xcvr._1_ ),
    .A2(net549),
    .B1(\u_usb_host.u_phy.usb_tx_dp_o ),
    .X(net83));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_usb_xcvr._6__549  (.HI(net549));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._7_  (.A(\u_usb_host.u_phy.usb_tx_oen_o ),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._8_  (.A(net44),
    .X(\u_usb_host.u_phy.usb_rx_dn_i ));
 sky130_fd_sc_hd__clkbuf_1 \u_usb_host.u_usb_xcvr._9_  (.A(net45),
    .X(\u_usb_host.u_phy.usb_rx_dp_i ));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_wb_rst._1_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net563),
    .RESET_B(net46),
    .Q(\u_usb_host.u_wb_rst.in_data_s ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_wb_rst._1__563  (.HI(net563));
 sky130_fd_sc_hd__dfrtp_1 \u_usb_host.u_wb_rst._2_  (.CLK(clknet_1_0__leaf_app_clk),
    .D(net659),
    .RESET_B(net46),
    .Q(\u_usb_host.u_wb_rst.in_data_2s ));
 sky130_fd_sc_hd__mux2_1 \u_usb_host.u_wb_rst.u_buf.genblk1.u_mux  (.A0(net570),
    .A1(net46),
    .S(net546),
    .X(\u_usb_host.u_async_wb.u_cmd_if.wr_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_usb_host.u_wb_rst.u_buf.genblk1.u_mux_546  (.LO(net546));
 sky130_fd_sc_hd__buf_4 wire2 (.A(net566),
    .X(net565));
 sky130_fd_sc_hd__clkbuf_2 wire3 (.A(usb_clk),
    .X(net566));
endmodule

