magic
tech sky130A
magscale 1 2
timestamp 1698826261
<< obsli1 >>
rect 1104 2159 18860 17425
<< obsm1 >>
rect 14 960 19950 17536
<< metal2 >>
rect 110 19200 166 20000
rect 294 19200 350 20000
rect 478 19200 534 20000
rect 662 19200 718 20000
rect 846 19200 902 20000
rect 1030 19200 1086 20000
rect 1214 19200 1270 20000
rect 1398 19200 1454 20000
rect 1582 19200 1638 20000
rect 1766 19200 1822 20000
rect 1950 19200 2006 20000
rect 2134 19200 2190 20000
rect 2318 19200 2374 20000
rect 110 0 166 800
rect 294 0 350 800
<< obsm2 >>
rect 18 19144 54 19200
rect 222 19144 238 19200
rect 406 19144 422 19200
rect 590 19144 606 19200
rect 774 19144 790 19200
rect 958 19144 974 19200
rect 1142 19144 1158 19200
rect 1326 19144 1342 19200
rect 1510 19144 1526 19200
rect 1694 19144 1710 19200
rect 1878 19144 1894 19200
rect 2062 19144 2078 19200
rect 2246 19144 2262 19200
rect 2430 19144 19944 19200
rect 18 856 19944 19144
rect 18 167 54 856
rect 222 167 238 856
rect 406 167 19944 856
<< metal3 >>
rect 0 4224 800 4344
rect 0 3952 800 4072
rect 0 3680 800 3800
rect 0 3408 800 3528
rect 0 3136 800 3256
rect 0 2864 800 2984
rect 0 2592 800 2712
rect 0 2320 800 2440
rect 0 2048 800 2168
rect 0 1776 800 1896
rect 0 1504 800 1624
rect 0 1232 800 1352
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
rect 19200 1504 20000 1624
rect 19200 1232 20000 1352
rect 19200 960 20000 1080
rect 19200 688 20000 808
rect 19200 416 20000 536
rect 19200 144 20000 264
<< obsm3 >>
rect 13 4424 19859 17441
rect 880 1704 19859 4424
rect 880 171 19120 1704
<< metal4 >>
rect 1484 2128 2724 17456
rect 5484 2128 6724 17456
rect 9484 2128 10724 17456
rect 13484 2128 14724 17456
rect 17484 2128 18724 17456
<< obsm4 >>
rect 18827 4115 19261 11661
<< labels >>
rlabel metal4 s 5484 2128 6724 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 13484 2128 14724 17456 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 1484 2128 2724 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 9484 2128 10724 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 17484 2128 18724 17456 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 0 416 800 536 6 clockp[0]
port 3 nsew signal output
rlabel metal3 s 0 144 800 264 6 clockp[1]
port 4 nsew signal output
rlabel metal3 s 0 2320 800 2440 6 dco
port 5 nsew signal input
rlabel metal3 s 0 1776 800 1896 6 div[0]
port 6 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 div[1]
port 7 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 div[2]
port 8 nsew signal input
rlabel metal3 s 0 960 800 1080 6 div[3]
port 9 nsew signal input
rlabel metal3 s 0 688 800 808 6 div[4]
port 10 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 enable
port 11 nsew signal input
rlabel metal3 s 0 4224 800 4344 6 ext_trim[0]
port 12 nsew signal input
rlabel metal2 s 2318 19200 2374 20000 6 ext_trim[10]
port 13 nsew signal input
rlabel metal2 s 2134 19200 2190 20000 6 ext_trim[11]
port 14 nsew signal input
rlabel metal2 s 1950 19200 2006 20000 6 ext_trim[12]
port 15 nsew signal input
rlabel metal2 s 1766 19200 1822 20000 6 ext_trim[13]
port 16 nsew signal input
rlabel metal2 s 1582 19200 1638 20000 6 ext_trim[14]
port 17 nsew signal input
rlabel metal2 s 1398 19200 1454 20000 6 ext_trim[15]
port 18 nsew signal input
rlabel metal2 s 1214 19200 1270 20000 6 ext_trim[16]
port 19 nsew signal input
rlabel metal2 s 1030 19200 1086 20000 6 ext_trim[17]
port 20 nsew signal input
rlabel metal2 s 846 19200 902 20000 6 ext_trim[18]
port 21 nsew signal input
rlabel metal2 s 662 19200 718 20000 6 ext_trim[19]
port 22 nsew signal input
rlabel metal3 s 0 3952 800 4072 6 ext_trim[1]
port 23 nsew signal input
rlabel metal3 s 19200 1504 20000 1624 6 ext_trim[20]
port 24 nsew signal input
rlabel metal3 s 19200 1232 20000 1352 6 ext_trim[21]
port 25 nsew signal input
rlabel metal3 s 19200 960 20000 1080 6 ext_trim[22]
port 26 nsew signal input
rlabel metal3 s 19200 688 20000 808 6 ext_trim[23]
port 27 nsew signal input
rlabel metal3 s 19200 416 20000 536 6 ext_trim[24]
port 28 nsew signal input
rlabel metal3 s 19200 144 20000 264 6 ext_trim[25]
port 29 nsew signal input
rlabel metal3 s 0 3680 800 3800 6 ext_trim[2]
port 30 nsew signal input
rlabel metal3 s 0 3408 800 3528 6 ext_trim[3]
port 31 nsew signal input
rlabel metal3 s 0 3136 800 3256 6 ext_trim[4]
port 32 nsew signal input
rlabel metal3 s 0 2864 800 2984 6 ext_trim[5]
port 33 nsew signal input
rlabel metal3 s 0 2592 800 2712 6 ext_trim[6]
port 34 nsew signal input
rlabel metal2 s 110 19200 166 20000 6 ext_trim[7]
port 35 nsew signal input
rlabel metal2 s 294 19200 350 20000 6 ext_trim[8]
port 36 nsew signal input
rlabel metal2 s 478 19200 534 20000 6 ext_trim[9]
port 37 nsew signal input
rlabel metal2 s 294 0 350 800 6 osc
port 38 nsew signal input
rlabel metal2 s 110 0 166 800 6 resetb
port 39 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 20000 20000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1608482
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/dg_pll/runs/dg_pll/results/signoff/dg_pll.magic.gds
string GDS_START 376646
<< end >>

