magic
tech sky130A
magscale 1 2
timestamp 1698751204
<< obsli1 >>
rect 1104 2159 98808 137649
<< obsm1 >>
rect 106 892 98808 138168
<< metal2 >>
rect 110 139200 166 140000
rect 294 139200 350 140000
rect 478 139200 534 140000
rect 662 139200 718 140000
rect 846 139200 902 140000
rect 1030 139200 1086 140000
rect 110 0 166 800
rect 294 0 350 800
<< obsm2 >>
rect 222 139144 238 139346
rect 406 139144 422 139346
rect 590 139144 606 139346
rect 774 139144 790 139346
rect 958 139144 974 139346
rect 1142 139144 94970 139346
rect 112 856 94970 139144
rect 222 800 238 856
rect 406 800 94970 856
<< metal3 >>
rect 0 101600 800 101720
rect 0 101328 800 101448
rect 0 101056 800 101176
rect 0 100784 800 100904
rect 0 100512 800 100632
rect 0 100240 800 100360
rect 0 99968 800 100088
rect 0 99696 800 99816
rect 0 99424 800 99544
rect 0 99152 800 99272
rect 0 98880 800 99000
rect 0 98608 800 98728
rect 0 98336 800 98456
rect 0 98064 800 98184
rect 0 97792 800 97912
rect 0 97520 800 97640
rect 0 97248 800 97368
rect 0 96976 800 97096
rect 0 96704 800 96824
rect 0 96432 800 96552
rect 0 96160 800 96280
rect 0 95888 800 96008
rect 0 95616 800 95736
rect 0 95344 800 95464
rect 0 95072 800 95192
rect 0 94800 800 94920
rect 0 94528 800 94648
rect 0 94256 800 94376
rect 0 93984 800 94104
rect 0 93712 800 93832
rect 0 93440 800 93560
rect 0 93168 800 93288
rect 0 92896 800 93016
rect 0 92624 800 92744
rect 0 92352 800 92472
rect 0 92080 800 92200
rect 0 91808 800 91928
rect 0 91536 800 91656
rect 0 91264 800 91384
rect 0 90992 800 91112
rect 0 90720 800 90840
rect 0 90448 800 90568
rect 0 90176 800 90296
rect 0 89904 800 90024
rect 0 89632 800 89752
rect 0 89360 800 89480
rect 0 89088 800 89208
rect 0 88816 800 88936
rect 0 88544 800 88664
rect 0 88272 800 88392
rect 0 88000 800 88120
rect 0 87728 800 87848
rect 0 87456 800 87576
rect 0 87184 800 87304
rect 0 86912 800 87032
rect 0 86640 800 86760
rect 0 86368 800 86488
rect 0 86096 800 86216
rect 0 85824 800 85944
rect 0 85552 800 85672
rect 0 85280 800 85400
rect 0 85008 800 85128
rect 0 84736 800 84856
rect 0 84464 800 84584
rect 0 84192 800 84312
rect 0 83920 800 84040
rect 0 83648 800 83768
rect 0 83376 800 83496
rect 0 83104 800 83224
rect 0 82832 800 82952
rect 0 82560 800 82680
rect 0 82288 800 82408
rect 0 82016 800 82136
rect 0 81744 800 81864
rect 0 81472 800 81592
rect 0 81200 800 81320
rect 0 80928 800 81048
rect 0 80656 800 80776
rect 0 80384 800 80504
rect 0 80112 800 80232
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
<< obsm3 >>
rect 800 101800 94966 137665
rect 880 80032 94966 101800
rect 800 61952 94966 80032
rect 880 60040 94966 61952
rect 800 2143 94966 60040
<< metal4 >>
rect 3748 2128 4988 137680
rect 13748 2128 14988 137680
rect 23748 2128 24988 137680
rect 33748 2128 34988 137680
rect 43748 2128 44988 137680
rect 53748 2128 54988 137680
rect 63748 2128 64988 137680
rect 73748 2128 74988 137680
rect 83748 2128 84988 137680
rect 93748 2128 94988 137680
<< obsm4 >>
rect 1899 27507 3668 133925
rect 5068 27507 13668 133925
rect 15068 27507 23668 133925
rect 25068 27507 33668 133925
rect 35068 27507 43668 133925
rect 45068 27507 53668 133925
rect 55068 27507 63668 133925
rect 65068 27507 65997 133925
<< labels >>
rlabel metal3 s 0 61752 800 61872 6 app_clk
port 1 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 cfg_cska_usb[0]
port 2 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 cfg_cska_usb[1]
port 3 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 cfg_cska_usb[2]
port 4 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 cfg_cska_usb[3]
port 5 nsew signal input
rlabel metal3 s 0 101600 800 101720 6 reg_ack
port 6 nsew signal output
rlabel metal3 s 0 82832 800 82952 6 reg_addr[0]
port 7 nsew signal input
rlabel metal3 s 0 82560 800 82680 6 reg_addr[1]
port 8 nsew signal input
rlabel metal3 s 0 82288 800 82408 6 reg_addr[2]
port 9 nsew signal input
rlabel metal3 s 0 82016 800 82136 6 reg_addr[3]
port 10 nsew signal input
rlabel metal3 s 0 81744 800 81864 6 reg_addr[4]
port 11 nsew signal input
rlabel metal3 s 0 81472 800 81592 6 reg_addr[5]
port 12 nsew signal input
rlabel metal3 s 0 81200 800 81320 6 reg_addr[6]
port 13 nsew signal input
rlabel metal3 s 0 80928 800 81048 6 reg_addr[7]
port 14 nsew signal input
rlabel metal3 s 0 80656 800 80776 6 reg_addr[8]
port 15 nsew signal input
rlabel metal3 s 0 83920 800 84040 6 reg_be[0]
port 16 nsew signal input
rlabel metal3 s 0 83648 800 83768 6 reg_be[1]
port 17 nsew signal input
rlabel metal3 s 0 83376 800 83496 6 reg_be[2]
port 18 nsew signal input
rlabel metal3 s 0 83104 800 83224 6 reg_be[3]
port 19 nsew signal input
rlabel metal3 s 0 80112 800 80232 6 reg_cs
port 20 nsew signal input
rlabel metal3 s 0 101328 800 101448 6 reg_rdata[0]
port 21 nsew signal output
rlabel metal3 s 0 98608 800 98728 6 reg_rdata[10]
port 22 nsew signal output
rlabel metal3 s 0 98336 800 98456 6 reg_rdata[11]
port 23 nsew signal output
rlabel metal3 s 0 98064 800 98184 6 reg_rdata[12]
port 24 nsew signal output
rlabel metal3 s 0 97792 800 97912 6 reg_rdata[13]
port 25 nsew signal output
rlabel metal3 s 0 97520 800 97640 6 reg_rdata[14]
port 26 nsew signal output
rlabel metal3 s 0 97248 800 97368 6 reg_rdata[15]
port 27 nsew signal output
rlabel metal3 s 0 96976 800 97096 6 reg_rdata[16]
port 28 nsew signal output
rlabel metal3 s 0 96704 800 96824 6 reg_rdata[17]
port 29 nsew signal output
rlabel metal3 s 0 96432 800 96552 6 reg_rdata[18]
port 30 nsew signal output
rlabel metal3 s 0 96160 800 96280 6 reg_rdata[19]
port 31 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 reg_rdata[1]
port 32 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 reg_rdata[20]
port 33 nsew signal output
rlabel metal3 s 0 95616 800 95736 6 reg_rdata[21]
port 34 nsew signal output
rlabel metal3 s 0 95344 800 95464 6 reg_rdata[22]
port 35 nsew signal output
rlabel metal3 s 0 95072 800 95192 6 reg_rdata[23]
port 36 nsew signal output
rlabel metal3 s 0 94800 800 94920 6 reg_rdata[24]
port 37 nsew signal output
rlabel metal3 s 0 94528 800 94648 6 reg_rdata[25]
port 38 nsew signal output
rlabel metal3 s 0 94256 800 94376 6 reg_rdata[26]
port 39 nsew signal output
rlabel metal3 s 0 93984 800 94104 6 reg_rdata[27]
port 40 nsew signal output
rlabel metal3 s 0 93712 800 93832 6 reg_rdata[28]
port 41 nsew signal output
rlabel metal3 s 0 93440 800 93560 6 reg_rdata[29]
port 42 nsew signal output
rlabel metal3 s 0 100784 800 100904 6 reg_rdata[2]
port 43 nsew signal output
rlabel metal3 s 0 93168 800 93288 6 reg_rdata[30]
port 44 nsew signal output
rlabel metal3 s 0 92896 800 93016 6 reg_rdata[31]
port 45 nsew signal output
rlabel metal3 s 0 100512 800 100632 6 reg_rdata[3]
port 46 nsew signal output
rlabel metal3 s 0 100240 800 100360 6 reg_rdata[4]
port 47 nsew signal output
rlabel metal3 s 0 99968 800 100088 6 reg_rdata[5]
port 48 nsew signal output
rlabel metal3 s 0 99696 800 99816 6 reg_rdata[6]
port 49 nsew signal output
rlabel metal3 s 0 99424 800 99544 6 reg_rdata[7]
port 50 nsew signal output
rlabel metal3 s 0 99152 800 99272 6 reg_rdata[8]
port 51 nsew signal output
rlabel metal3 s 0 98880 800 99000 6 reg_rdata[9]
port 52 nsew signal output
rlabel metal3 s 0 92624 800 92744 6 reg_wdata[0]
port 53 nsew signal input
rlabel metal3 s 0 89904 800 90024 6 reg_wdata[10]
port 54 nsew signal input
rlabel metal3 s 0 89632 800 89752 6 reg_wdata[11]
port 55 nsew signal input
rlabel metal3 s 0 89360 800 89480 6 reg_wdata[12]
port 56 nsew signal input
rlabel metal3 s 0 89088 800 89208 6 reg_wdata[13]
port 57 nsew signal input
rlabel metal3 s 0 88816 800 88936 6 reg_wdata[14]
port 58 nsew signal input
rlabel metal3 s 0 88544 800 88664 6 reg_wdata[15]
port 59 nsew signal input
rlabel metal3 s 0 88272 800 88392 6 reg_wdata[16]
port 60 nsew signal input
rlabel metal3 s 0 88000 800 88120 6 reg_wdata[17]
port 61 nsew signal input
rlabel metal3 s 0 87728 800 87848 6 reg_wdata[18]
port 62 nsew signal input
rlabel metal3 s 0 87456 800 87576 6 reg_wdata[19]
port 63 nsew signal input
rlabel metal3 s 0 92352 800 92472 6 reg_wdata[1]
port 64 nsew signal input
rlabel metal3 s 0 87184 800 87304 6 reg_wdata[20]
port 65 nsew signal input
rlabel metal3 s 0 86912 800 87032 6 reg_wdata[21]
port 66 nsew signal input
rlabel metal3 s 0 86640 800 86760 6 reg_wdata[22]
port 67 nsew signal input
rlabel metal3 s 0 86368 800 86488 6 reg_wdata[23]
port 68 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 reg_wdata[24]
port 69 nsew signal input
rlabel metal3 s 0 85824 800 85944 6 reg_wdata[25]
port 70 nsew signal input
rlabel metal3 s 0 85552 800 85672 6 reg_wdata[26]
port 71 nsew signal input
rlabel metal3 s 0 85280 800 85400 6 reg_wdata[27]
port 72 nsew signal input
rlabel metal3 s 0 85008 800 85128 6 reg_wdata[28]
port 73 nsew signal input
rlabel metal3 s 0 84736 800 84856 6 reg_wdata[29]
port 74 nsew signal input
rlabel metal3 s 0 92080 800 92200 6 reg_wdata[2]
port 75 nsew signal input
rlabel metal3 s 0 84464 800 84584 6 reg_wdata[30]
port 76 nsew signal input
rlabel metal3 s 0 84192 800 84312 6 reg_wdata[31]
port 77 nsew signal input
rlabel metal3 s 0 91808 800 91928 6 reg_wdata[3]
port 78 nsew signal input
rlabel metal3 s 0 91536 800 91656 6 reg_wdata[4]
port 79 nsew signal input
rlabel metal3 s 0 91264 800 91384 6 reg_wdata[5]
port 80 nsew signal input
rlabel metal3 s 0 90992 800 91112 6 reg_wdata[6]
port 81 nsew signal input
rlabel metal3 s 0 90720 800 90840 6 reg_wdata[7]
port 82 nsew signal input
rlabel metal3 s 0 90448 800 90568 6 reg_wdata[8]
port 83 nsew signal input
rlabel metal3 s 0 90176 800 90296 6 reg_wdata[9]
port 84 nsew signal input
rlabel metal3 s 0 80384 800 80504 6 reg_wr
port 85 nsew signal input
rlabel metal2 s 110 0 166 800 6 usb_clk
port 86 nsew signal input
rlabel metal2 s 294 139200 350 140000 6 usb_in_dn
port 87 nsew signal input
rlabel metal2 s 110 139200 166 140000 6 usb_in_dp
port 88 nsew signal input
rlabel metal2 s 1030 139200 1086 140000 6 usb_intr_o
port 89 nsew signal output
rlabel metal2 s 662 139200 718 140000 6 usb_out_dn
port 90 nsew signal output
rlabel metal2 s 478 139200 534 140000 6 usb_out_dp
port 91 nsew signal output
rlabel metal2 s 846 139200 902 140000 6 usb_out_tx_oen
port 92 nsew signal output
rlabel metal2 s 294 0 350 800 6 usb_rstn
port 93 nsew signal input
rlabel metal4 s 3748 2128 4988 137680 6 vccd1
port 94 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 137680 6 vccd1
port 94 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 137680 6 vccd1
port 94 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 137680 6 vccd1
port 94 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 137680 6 vccd1
port 94 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 137680 6 vssd1
port 95 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 137680 6 vssd1
port 95 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 137680 6 vssd1
port 95 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 137680 6 vssd1
port 95 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 137680 6 vssd1
port 95 nsew ground bidirectional
rlabel metal3 s 0 61208 800 61328 6 wbd_clk_int
port 96 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 wbd_clk_usb
port 97 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100000 140000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22840512
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/usb_top/runs/usb_top/results/signoff/usb_top.magic.gds
string GDS_START 947178
<< end >>

