VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO bus_rep_south
  CLASS BLOCK ;
  FOREIGN bus_rep_south ;
  ORIGIN 0.000 0.000 ;
  SIZE 2650.000 BY 60.000 ;
  PIN ch_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 0.370 0.000 0.650 4.000 ;
    END
  END ch_in[0]
  PIN ch_in[100]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 544.370 0.000 544.650 4.000 ;
    END
  END ch_in[100]
  PIN ch_in[101]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 549.810 0.000 550.090 4.000 ;
    END
  END ch_in[101]
  PIN ch_in[102]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1277.750 56.000 1278.030 60.000 ;
    END
  END ch_in[102]
  PIN ch_in[103]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 560.690 0.000 560.970 4.000 ;
    END
  END ch_in[103]
  PIN ch_in[104]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 566.130 0.000 566.410 4.000 ;
    END
  END ch_in[104]
  PIN ch_in[105]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1285.910 56.000 1286.190 60.000 ;
    END
  END ch_in[105]
  PIN ch_in[106]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 600.130 0.000 600.410 4.000 ;
    END
  END ch_in[106]
  PIN ch_in[107]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1803.050 56.000 1803.330 60.000 ;
    END
  END ch_in[107]
  PIN ch_in[108]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 621.890 0.000 622.170 4.000 ;
    END
  END ch_in[108]
  PIN ch_in[109]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1808.490 56.000 1808.770 60.000 ;
    END
  END ch_in[109]
  PIN ch_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 54.770 0.000 55.050 4.000 ;
    END
  END ch_in[10]
  PIN ch_in[110]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 643.650 0.000 643.930 4.000 ;
    END
  END ch_in[110]
  PIN ch_in[111]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1813.930 56.000 1814.210 60.000 ;
    END
  END ch_in[111]
  PIN ch_in[112]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 665.410 0.000 665.690 4.000 ;
    END
  END ch_in[112]
  PIN ch_in[113]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1819.370 56.000 1819.650 60.000 ;
    END
  END ch_in[113]
  PIN ch_in[114]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 687.170 0.000 687.450 4.000 ;
    END
  END ch_in[114]
  PIN ch_in[115]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1824.810 56.000 1825.090 60.000 ;
    END
  END ch_in[115]
  PIN ch_in[116]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 708.930 0.000 709.210 4.000 ;
    END
  END ch_in[116]
  PIN ch_in[117]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1830.250 56.000 1830.530 60.000 ;
    END
  END ch_in[117]
  PIN ch_in[118]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 730.690 0.000 730.970 4.000 ;
    END
  END ch_in[118]
  PIN ch_in[119]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1835.690 56.000 1835.970 60.000 ;
    END
  END ch_in[119]
  PIN ch_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 60.210 0.000 60.490 4.000 ;
    END
  END ch_in[11]
  PIN ch_in[120]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 752.450 0.000 752.730 4.000 ;
    END
  END ch_in[120]
  PIN ch_in[121]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1841.130 56.000 1841.410 60.000 ;
    END
  END ch_in[121]
  PIN ch_in[122]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 774.210 0.000 774.490 4.000 ;
    END
  END ch_in[122]
  PIN ch_in[123]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1846.570 56.000 1846.850 60.000 ;
    END
  END ch_in[123]
  PIN ch_in[124]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 795.970 0.000 796.250 4.000 ;
    END
  END ch_in[124]
  PIN ch_in[125]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1852.010 56.000 1852.290 60.000 ;
    END
  END ch_in[125]
  PIN ch_in[126]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 810.250 0.000 810.530 4.000 ;
    END
  END ch_in[126]
  PIN ch_in[127]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1857.450 56.000 1857.730 60.000 ;
    END
  END ch_in[127]
  PIN ch_in[128]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 832.010 0.000 832.290 4.000 ;
    END
  END ch_in[128]
  PIN ch_in[129]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1862.890 56.000 1863.170 60.000 ;
    END
  END ch_in[129]
  PIN ch_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1032.950 56.000 1033.230 60.000 ;
    END
  END ch_in[12]
  PIN ch_in[130]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 853.770 0.000 854.050 4.000 ;
    END
  END ch_in[130]
  PIN ch_in[131]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1868.330 56.000 1868.610 60.000 ;
    END
  END ch_in[131]
  PIN ch_in[132]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 875.530 0.000 875.810 4.000 ;
    END
  END ch_in[132]
  PIN ch_in[133]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1873.770 56.000 1874.050 60.000 ;
    END
  END ch_in[133]
  PIN ch_in[134]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 897.290 0.000 897.570 4.000 ;
    END
  END ch_in[134]
  PIN ch_in[135]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1879.210 56.000 1879.490 60.000 ;
    END
  END ch_in[135]
  PIN ch_in[136]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 919.050 0.000 919.330 4.000 ;
    END
  END ch_in[136]
  PIN ch_in[137]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1884.650 56.000 1884.930 60.000 ;
    END
  END ch_in[137]
  PIN ch_in[138]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 940.810 0.000 941.090 4.000 ;
    END
  END ch_in[138]
  PIN ch_in[139]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1890.090 56.000 1890.370 60.000 ;
    END
  END ch_in[139]
  PIN ch_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 71.090 0.000 71.370 4.000 ;
    END
  END ch_in[13]
  PIN ch_in[140]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 962.570 0.000 962.850 4.000 ;
    END
  END ch_in[140]
  PIN ch_in[141]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1895.530 56.000 1895.810 60.000 ;
    END
  END ch_in[141]
  PIN ch_in[142]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1898.250 56.000 1898.530 60.000 ;
    END
  END ch_in[142]
  PIN ch_in[143]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1900.970 56.000 1901.250 60.000 ;
    END
  END ch_in[143]
  PIN ch_in[144]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1903.690 56.000 1903.970 60.000 ;
    END
  END ch_in[144]
  PIN ch_in[145]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1906.410 56.000 1906.690 60.000 ;
    END
  END ch_in[145]
  PIN ch_in[146]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1909.130 56.000 1909.410 60.000 ;
    END
  END ch_in[146]
  PIN ch_in[147]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1911.850 56.000 1912.130 60.000 ;
    END
  END ch_in[147]
  PIN ch_in[148]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1914.570 56.000 1914.850 60.000 ;
    END
  END ch_in[148]
  PIN ch_in[149]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1917.290 56.000 1917.570 60.000 ;
    END
  END ch_in[149]
  PIN ch_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 76.530 0.000 76.810 4.000 ;
    END
  END ch_in[14]
  PIN ch_in[150]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1920.010 56.000 1920.290 60.000 ;
    END
  END ch_in[150]
  PIN ch_in[151]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1922.730 55.860 1923.010 60.000 ;
    END
  END ch_in[151]
  PIN ch_in[152]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1925.450 56.000 1925.730 60.000 ;
    END
  END ch_in[152]
  PIN ch_in[153]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1928.170 56.000 1928.450 60.000 ;
    END
  END ch_in[153]
  PIN ch_in[154]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1930.890 56.000 1931.170 60.000 ;
    END
  END ch_in[154]
  PIN ch_in[155]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1933.610 56.000 1933.890 60.000 ;
    END
  END ch_in[155]
  PIN ch_in[156]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1936.330 56.000 1936.610 60.000 ;
    END
  END ch_in[156]
  PIN ch_in[157]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1939.050 56.000 1939.330 60.000 ;
    END
  END ch_in[157]
  PIN ch_in[158]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1941.770 56.000 1942.050 60.000 ;
    END
  END ch_in[158]
  PIN ch_in[159]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1944.490 56.000 1944.770 60.000 ;
    END
  END ch_in[159]
  PIN ch_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 81.970 0.000 82.250 4.000 ;
    END
  END ch_in[15]
  PIN ch_in[160]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1947.210 56.000 1947.490 60.000 ;
    END
  END ch_in[160]
  PIN ch_in[161]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1949.930 56.000 1950.210 60.000 ;
    END
  END ch_in[161]
  PIN ch_in[162]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1952.650 56.000 1952.930 60.000 ;
    END
  END ch_in[162]
  PIN ch_in[163]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1955.370 56.000 1955.650 60.000 ;
    END
  END ch_in[163]
  PIN ch_in[164]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1958.090 56.000 1958.370 60.000 ;
    END
  END ch_in[164]
  PIN ch_in[165]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1960.810 56.000 1961.090 60.000 ;
    END
  END ch_in[165]
  PIN ch_in[166]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1963.530 56.000 1963.810 60.000 ;
    END
  END ch_in[166]
  PIN ch_in[167]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1966.250 56.000 1966.530 60.000 ;
    END
  END ch_in[167]
  PIN ch_in[168]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1968.970 56.000 1969.250 60.000 ;
    END
  END ch_in[168]
  PIN ch_in[169]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1971.690 56.000 1971.970 60.000 ;
    END
  END ch_in[169]
  PIN ch_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1043.830 56.000 1044.110 60.000 ;
    END
  END ch_in[16]
  PIN ch_in[170]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1974.410 56.000 1974.690 60.000 ;
    END
  END ch_in[170]
  PIN ch_in[171]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1977.130 56.000 1977.410 60.000 ;
    END
  END ch_in[171]
  PIN ch_in[172]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1979.850 56.000 1980.130 60.000 ;
    END
  END ch_in[172]
  PIN ch_in[173]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1982.570 56.000 1982.850 60.000 ;
    END
  END ch_in[173]
  PIN ch_in[174]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1985.290 55.860 1985.570 60.000 ;
    END
  END ch_in[174]
  PIN ch_in[175]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1988.010 56.000 1988.290 60.000 ;
    END
  END ch_in[175]
  PIN ch_in[176]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1990.730 56.000 1991.010 60.000 ;
    END
  END ch_in[176]
  PIN ch_in[177]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1993.450 56.000 1993.730 60.000 ;
    END
  END ch_in[177]
  PIN ch_in[178]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1996.170 56.000 1996.450 60.000 ;
    END
  END ch_in[178]
  PIN ch_in[179]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1998.890 56.000 1999.170 60.000 ;
    END
  END ch_in[179]
  PIN ch_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 92.850 0.000 93.130 4.000 ;
    END
  END ch_in[17]
  PIN ch_in[180]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2001.610 56.000 2001.890 60.000 ;
    END
  END ch_in[180]
  PIN ch_in[181]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2004.330 56.000 2004.610 60.000 ;
    END
  END ch_in[181]
  PIN ch_in[182]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2007.050 56.000 2007.330 60.000 ;
    END
  END ch_in[182]
  PIN ch_in[183]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2009.770 56.000 2010.050 60.000 ;
    END
  END ch_in[183]
  PIN ch_in[184]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2012.490 56.000 2012.770 60.000 ;
    END
  END ch_in[184]
  PIN ch_in[185]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2015.210 56.000 2015.490 60.000 ;
    END
  END ch_in[185]
  PIN ch_in[186]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2017.930 56.000 2018.210 60.000 ;
    END
  END ch_in[186]
  PIN ch_in[187]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2020.650 56.000 2020.930 60.000 ;
    END
  END ch_in[187]
  PIN ch_in[188]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2200.170 56.000 2200.450 60.000 ;
    END
  END ch_in[188]
  PIN ch_in[189]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2201.530 56.000 2201.810 60.000 ;
    END
  END ch_in[189]
  PIN ch_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 98.290 0.000 98.570 4.000 ;
    END
  END ch_in[18]
  PIN ch_in[190]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2202.890 56.000 2203.170 60.000 ;
    END
  END ch_in[190]
  PIN ch_in[191]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2204.250 56.000 2204.530 60.000 ;
    END
  END ch_in[191]
  PIN ch_in[192]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2205.610 56.000 2205.890 60.000 ;
    END
  END ch_in[192]
  PIN ch_in[193]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2206.970 56.000 2207.250 60.000 ;
    END
  END ch_in[193]
  PIN ch_in[194]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2208.330 56.000 2208.610 60.000 ;
    END
  END ch_in[194]
  PIN ch_in[195]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2209.690 56.000 2209.970 60.000 ;
    END
  END ch_in[195]
  PIN ch_in[196]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2211.050 56.000 2211.330 60.000 ;
    END
  END ch_in[196]
  PIN ch_in[197]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2212.410 56.000 2212.690 60.000 ;
    END
  END ch_in[197]
  PIN ch_in[198]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2213.770 55.860 2214.050 60.000 ;
    END
  END ch_in[198]
  PIN ch_in[199]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2215.130 56.000 2215.410 60.000 ;
    END
  END ch_in[199]
  PIN ch_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 103.730 0.000 104.010 4.000 ;
    END
  END ch_in[19]
  PIN ch_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 5.810 0.000 6.090 4.000 ;
    END
  END ch_in[1]
  PIN ch_in[200]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2216.490 56.000 2216.770 60.000 ;
    END
  END ch_in[200]
  PIN ch_in[201]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2217.850 56.000 2218.130 60.000 ;
    END
  END ch_in[201]
  PIN ch_in[202]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2219.210 56.000 2219.490 60.000 ;
    END
  END ch_in[202]
  PIN ch_in[203]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2220.570 56.000 2220.850 60.000 ;
    END
  END ch_in[203]
  PIN ch_in[204]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2221.930 56.000 2222.210 60.000 ;
    END
  END ch_in[204]
  PIN ch_in[205]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2223.290 56.000 2223.570 60.000 ;
    END
  END ch_in[205]
  PIN ch_in[206]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2224.650 56.000 2224.930 60.000 ;
    END
  END ch_in[206]
  PIN ch_in[207]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2226.010 56.000 2226.290 60.000 ;
    END
  END ch_in[207]
  PIN ch_in[208]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2227.370 56.000 2227.650 60.000 ;
    END
  END ch_in[208]
  PIN ch_in[209]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2228.730 56.000 2229.010 60.000 ;
    END
  END ch_in[209]
  PIN ch_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1054.710 56.000 1054.990 60.000 ;
    END
  END ch_in[20]
  PIN ch_in[210]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2230.090 56.000 2230.370 60.000 ;
    END
  END ch_in[210]
  PIN ch_in[211]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2231.450 56.000 2231.730 60.000 ;
    END
  END ch_in[211]
  PIN ch_in[212]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2232.810 56.000 2233.090 60.000 ;
    END
  END ch_in[212]
  PIN ch_in[213]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2234.170 56.000 2234.450 60.000 ;
    END
  END ch_in[213]
  PIN ch_in[214]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2235.530 55.860 2235.810 60.000 ;
    END
  END ch_in[214]
  PIN ch_in[215]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2236.890 56.000 2237.170 60.000 ;
    END
  END ch_in[215]
  PIN ch_in[216]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2238.250 56.000 2238.530 60.000 ;
    END
  END ch_in[216]
  PIN ch_in[217]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2239.610 56.000 2239.890 60.000 ;
    END
  END ch_in[217]
  PIN ch_in[218]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2240.970 56.000 2241.250 60.000 ;
    END
  END ch_in[218]
  PIN ch_in[219]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2242.330 56.000 2242.610 60.000 ;
    END
  END ch_in[219]
  PIN ch_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 114.610 0.000 114.890 4.000 ;
    END
  END ch_in[21]
  PIN ch_in[220]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2400.090 56.000 2400.370 60.000 ;
    END
  END ch_in[220]
  PIN ch_in[221]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2401.450 55.860 2401.730 60.000 ;
    END
  END ch_in[221]
  PIN ch_in[222]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2402.810 56.000 2403.090 60.000 ;
    END
  END ch_in[222]
  PIN ch_in[223]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2404.170 56.000 2404.450 60.000 ;
    END
  END ch_in[223]
  PIN ch_in[224]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2405.530 56.000 2405.810 60.000 ;
    END
  END ch_in[224]
  PIN ch_in[225]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2406.890 56.000 2407.170 60.000 ;
    END
  END ch_in[225]
  PIN ch_in[226]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2408.250 56.000 2408.530 60.000 ;
    END
  END ch_in[226]
  PIN ch_in[227]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2409.610 56.000 2409.890 60.000 ;
    END
  END ch_in[227]
  PIN ch_in[228]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2410.970 56.000 2411.250 60.000 ;
    END
  END ch_in[228]
  PIN ch_in[229]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2412.330 56.000 2412.610 60.000 ;
    END
  END ch_in[229]
  PIN ch_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 120.050 0.000 120.330 4.000 ;
    END
  END ch_in[22]
  PIN ch_in[230]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2413.690 56.000 2413.970 60.000 ;
    END
  END ch_in[230]
  PIN ch_in[231]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2415.050 55.860 2415.330 60.000 ;
    END
  END ch_in[231]
  PIN ch_in[232]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2416.410 56.000 2416.690 60.000 ;
    END
  END ch_in[232]
  PIN ch_in[233]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2417.770 56.000 2418.050 60.000 ;
    END
  END ch_in[233]
  PIN ch_in[234]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2419.130 56.000 2419.410 60.000 ;
    END
  END ch_in[234]
  PIN ch_in[235]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2420.490 56.000 2420.770 60.000 ;
    END
  END ch_in[235]
  PIN ch_in[236]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2421.850 56.000 2422.130 60.000 ;
    END
  END ch_in[236]
  PIN ch_in[237]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2423.210 56.000 2423.490 60.000 ;
    END
  END ch_in[237]
  PIN ch_in[238]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2424.570 56.000 2424.850 60.000 ;
    END
  END ch_in[238]
  PIN ch_in[239]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2425.930 56.000 2426.210 60.000 ;
    END
  END ch_in[239]
  PIN ch_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 125.490 0.000 125.770 4.000 ;
    END
  END ch_in[23]
  PIN ch_in[240]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2427.290 56.000 2427.570 60.000 ;
    END
  END ch_in[240]
  PIN ch_in[241]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2428.650 56.000 2428.930 60.000 ;
    END
  END ch_in[241]
  PIN ch_in[242]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2430.010 56.000 2430.290 60.000 ;
    END
  END ch_in[242]
  PIN ch_in[243]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2431.370 56.000 2431.650 60.000 ;
    END
  END ch_in[243]
  PIN ch_in[244]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2432.730 56.000 2433.010 60.000 ;
    END
  END ch_in[244]
  PIN ch_in[245]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2434.090 56.000 2434.370 60.000 ;
    END
  END ch_in[245]
  PIN ch_in[246]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2435.450 56.000 2435.730 60.000 ;
    END
  END ch_in[246]
  PIN ch_in[247]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2436.810 56.000 2437.090 60.000 ;
    END
  END ch_in[247]
  PIN ch_in[248]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2438.170 56.000 2438.450 60.000 ;
    END
  END ch_in[248]
  PIN ch_in[249]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2439.530 56.000 2439.810 60.000 ;
    END
  END ch_in[249]
  PIN ch_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1065.590 56.000 1065.870 60.000 ;
    END
  END ch_in[24]
  PIN ch_in[250]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2440.890 56.000 2441.170 60.000 ;
    END
  END ch_in[250]
  PIN ch_in[251]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2442.250 56.000 2442.530 60.000 ;
    END
  END ch_in[251]
  PIN ch_in[252]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2496.650 0.000 2496.930 4.000 ;
    END
  END ch_in[252]
  PIN ch_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 136.370 0.000 136.650 4.000 ;
    END
  END ch_in[25]
  PIN ch_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 141.810 0.000 142.090 4.000 ;
    END
  END ch_in[26]
  PIN ch_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1073.750 56.000 1074.030 60.000 ;
    END
  END ch_in[27]
  PIN ch_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 152.690 0.000 152.970 4.000 ;
    END
  END ch_in[28]
  PIN ch_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 158.130 0.000 158.410 4.000 ;
    END
  END ch_in[29]
  PIN ch_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1005.750 56.000 1006.030 60.000 ;
    END
  END ch_in[2]
  PIN ch_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1081.910 56.000 1082.190 60.000 ;
    END
  END ch_in[30]
  PIN ch_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 169.010 0.000 169.290 4.000 ;
    END
  END ch_in[31]
  PIN ch_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 174.450 0.000 174.730 4.000 ;
    END
  END ch_in[32]
  PIN ch_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1090.070 56.000 1090.350 60.000 ;
    END
  END ch_in[33]
  PIN ch_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 185.330 0.000 185.610 4.000 ;
    END
  END ch_in[34]
  PIN ch_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 190.770 0.000 191.050 4.000 ;
    END
  END ch_in[35]
  PIN ch_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1098.230 56.000 1098.510 60.000 ;
    END
  END ch_in[36]
  PIN ch_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 201.650 0.000 201.930 4.000 ;
    END
  END ch_in[37]
  PIN ch_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 207.090 0.000 207.370 4.000 ;
    END
  END ch_in[38]
  PIN ch_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1106.390 56.000 1106.670 60.000 ;
    END
  END ch_in[39]
  PIN ch_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 16.690 0.000 16.970 4.000 ;
    END
  END ch_in[3]
  PIN ch_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 217.970 0.000 218.250 4.000 ;
    END
  END ch_in[40]
  PIN ch_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 223.410 0.000 223.690 4.000 ;
    END
  END ch_in[41]
  PIN ch_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1114.550 56.000 1114.830 60.000 ;
    END
  END ch_in[42]
  PIN ch_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 234.290 0.000 234.570 4.000 ;
    END
  END ch_in[43]
  PIN ch_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 239.730 0.000 240.010 4.000 ;
    END
  END ch_in[44]
  PIN ch_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1122.710 56.000 1122.990 60.000 ;
    END
  END ch_in[45]
  PIN ch_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 250.610 0.000 250.890 4.000 ;
    END
  END ch_in[46]
  PIN ch_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 256.050 0.000 256.330 4.000 ;
    END
  END ch_in[47]
  PIN ch_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1130.870 56.000 1131.150 60.000 ;
    END
  END ch_in[48]
  PIN ch_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 266.930 0.000 267.210 4.000 ;
    END
  END ch_in[49]
  PIN ch_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 22.130 0.000 22.410 4.000 ;
    END
  END ch_in[4]
  PIN ch_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 272.370 0.000 272.650 4.000 ;
    END
  END ch_in[50]
  PIN ch_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1139.030 56.000 1139.310 60.000 ;
    END
  END ch_in[51]
  PIN ch_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 283.250 0.000 283.530 4.000 ;
    END
  END ch_in[52]
  PIN ch_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 288.690 0.000 288.970 4.000 ;
    END
  END ch_in[53]
  PIN ch_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1147.190 56.000 1147.470 60.000 ;
    END
  END ch_in[54]
  PIN ch_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 299.570 0.000 299.850 4.000 ;
    END
  END ch_in[55]
  PIN ch_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 305.010 0.000 305.290 4.000 ;
    END
  END ch_in[56]
  PIN ch_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1155.350 56.000 1155.630 60.000 ;
    END
  END ch_in[57]
  PIN ch_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 315.890 0.000 316.170 4.000 ;
    END
  END ch_in[58]
  PIN ch_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 321.330 0.000 321.610 4.000 ;
    END
  END ch_in[59]
  PIN ch_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 27.570 0.000 27.850 4.000 ;
    END
  END ch_in[5]
  PIN ch_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1163.510 56.000 1163.790 60.000 ;
    END
  END ch_in[60]
  PIN ch_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END ch_in[61]
  PIN ch_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 337.650 0.000 337.930 4.000 ;
    END
  END ch_in[62]
  PIN ch_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1171.670 56.000 1171.950 60.000 ;
    END
  END ch_in[63]
  PIN ch_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 348.530 0.000 348.810 4.000 ;
    END
  END ch_in[64]
  PIN ch_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 353.970 0.000 354.250 4.000 ;
    END
  END ch_in[65]
  PIN ch_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1179.830 56.000 1180.110 60.000 ;
    END
  END ch_in[66]
  PIN ch_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 364.850 0.000 365.130 4.000 ;
    END
  END ch_in[67]
  PIN ch_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 370.290 0.000 370.570 4.000 ;
    END
  END ch_in[68]
  PIN ch_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1187.990 56.000 1188.270 60.000 ;
    END
  END ch_in[69]
  PIN ch_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 33.010 0.000 33.290 4.000 ;
    END
  END ch_in[6]
  PIN ch_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 381.170 0.000 381.450 4.000 ;
    END
  END ch_in[70]
  PIN ch_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 386.610 0.000 386.890 4.000 ;
    END
  END ch_in[71]
  PIN ch_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1196.150 56.000 1196.430 60.000 ;
    END
  END ch_in[72]
  PIN ch_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 397.490 0.000 397.770 4.000 ;
    END
  END ch_in[73]
  PIN ch_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 402.930 0.000 403.210 4.000 ;
    END
  END ch_in[74]
  PIN ch_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1204.310 56.000 1204.590 60.000 ;
    END
  END ch_in[75]
  PIN ch_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 413.810 0.000 414.090 4.000 ;
    END
  END ch_in[76]
  PIN ch_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 419.250 0.000 419.530 4.000 ;
    END
  END ch_in[77]
  PIN ch_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1212.470 56.000 1212.750 60.000 ;
    END
  END ch_in[78]
  PIN ch_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 430.130 0.000 430.410 4.000 ;
    END
  END ch_in[79]
  PIN ch_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 38.450 0.000 38.730 4.000 ;
    END
  END ch_in[7]
  PIN ch_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 435.570 0.000 435.850 4.000 ;
    END
  END ch_in[80]
  PIN ch_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1220.630 55.860 1220.910 60.000 ;
    END
  END ch_in[81]
  PIN ch_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 446.450 0.000 446.730 4.000 ;
    END
  END ch_in[82]
  PIN ch_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 451.890 0.000 452.170 4.000 ;
    END
  END ch_in[83]
  PIN ch_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1228.790 56.000 1229.070 60.000 ;
    END
  END ch_in[84]
  PIN ch_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 462.770 0.000 463.050 4.000 ;
    END
  END ch_in[85]
  PIN ch_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 468.210 0.000 468.490 4.000 ;
    END
  END ch_in[86]
  PIN ch_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1236.950 56.000 1237.230 60.000 ;
    END
  END ch_in[87]
  PIN ch_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 479.090 0.000 479.370 4.000 ;
    END
  END ch_in[88]
  PIN ch_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 484.530 0.000 484.810 4.000 ;
    END
  END ch_in[89]
  PIN ch_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1022.070 56.000 1022.350 60.000 ;
    END
  END ch_in[8]
  PIN ch_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1245.110 56.000 1245.390 60.000 ;
    END
  END ch_in[90]
  PIN ch_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 495.410 0.000 495.690 4.000 ;
    END
  END ch_in[91]
  PIN ch_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 500.850 0.000 501.130 4.000 ;
    END
  END ch_in[92]
  PIN ch_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1253.270 56.000 1253.550 60.000 ;
    END
  END ch_in[93]
  PIN ch_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 511.730 0.000 512.010 4.000 ;
    END
  END ch_in[94]
  PIN ch_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 517.170 0.000 517.450 4.000 ;
    END
  END ch_in[95]
  PIN ch_in[96]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1261.430 56.000 1261.710 60.000 ;
    END
  END ch_in[96]
  PIN ch_in[97]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 528.050 0.000 528.330 4.000 ;
    END
  END ch_in[97]
  PIN ch_in[98]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 533.490 0.000 533.770 4.000 ;
    END
  END ch_in[98]
  PIN ch_in[99]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1269.590 56.000 1269.870 60.000 ;
    END
  END ch_in[99]
  PIN ch_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 49.330 0.000 49.610 4.000 ;
    END
  END ch_in[9]
  PIN ch_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1000.310 56.000 1000.590 60.000 ;
    END
  END ch_out[0]
  PIN ch_out[100]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1272.310 56.000 1272.590 60.000 ;
    END
  END ch_out[100]
  PIN ch_out[101]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1275.030 56.000 1275.310 60.000 ;
    END
  END ch_out[101]
  PIN ch_out[102]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 555.250 0.000 555.530 4.000 ;
    END
  END ch_out[102]
  PIN ch_out[103]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1280.470 56.000 1280.750 60.000 ;
    END
  END ch_out[103]
  PIN ch_out[104]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1283.190 56.000 1283.470 60.000 ;
    END
  END ch_out[104]
  PIN ch_out[105]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 571.570 0.000 571.850 4.000 ;
    END
  END ch_out[105]
  PIN ch_out[106]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1800.330 56.000 1800.610 60.000 ;
    END
  END ch_out[106]
  PIN ch_out[107]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 611.010 0.000 611.290 4.000 ;
    END
  END ch_out[107]
  PIN ch_out[108]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1805.770 56.000 1806.050 60.000 ;
    END
  END ch_out[108]
  PIN ch_out[109]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 632.770 0.000 633.050 4.000 ;
    END
  END ch_out[109]
  PIN ch_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1027.510 56.000 1027.790 60.000 ;
    END
  END ch_out[10]
  PIN ch_out[110]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1811.210 56.000 1811.490 60.000 ;
    END
  END ch_out[110]
  PIN ch_out[111]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 654.530 0.000 654.810 4.000 ;
    END
  END ch_out[111]
  PIN ch_out[112]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1816.650 56.000 1816.930 60.000 ;
    END
  END ch_out[112]
  PIN ch_out[113]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 676.290 0.000 676.570 4.000 ;
    END
  END ch_out[113]
  PIN ch_out[114]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1822.090 56.000 1822.370 60.000 ;
    END
  END ch_out[114]
  PIN ch_out[115]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 698.050 0.000 698.330 4.000 ;
    END
  END ch_out[115]
  PIN ch_out[116]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1827.530 56.000 1827.810 60.000 ;
    END
  END ch_out[116]
  PIN ch_out[117]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 719.810 0.000 720.090 4.000 ;
    END
  END ch_out[117]
  PIN ch_out[118]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1832.970 56.000 1833.250 60.000 ;
    END
  END ch_out[118]
  PIN ch_out[119]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 741.570 0.000 741.850 4.000 ;
    END
  END ch_out[119]
  PIN ch_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1030.230 56.000 1030.510 60.000 ;
    END
  END ch_out[11]
  PIN ch_out[120]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1838.410 56.000 1838.690 60.000 ;
    END
  END ch_out[120]
  PIN ch_out[121]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 763.330 0.000 763.610 4.000 ;
    END
  END ch_out[121]
  PIN ch_out[122]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1843.850 56.000 1844.130 60.000 ;
    END
  END ch_out[122]
  PIN ch_out[123]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 785.090 0.000 785.370 4.000 ;
    END
  END ch_out[123]
  PIN ch_out[124]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1849.290 56.000 1849.570 60.000 ;
    END
  END ch_out[124]
  PIN ch_out[125]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 806.850 0.000 807.130 4.000 ;
    END
  END ch_out[125]
  PIN ch_out[126]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1854.730 56.000 1855.010 60.000 ;
    END
  END ch_out[126]
  PIN ch_out[127]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 821.130 0.000 821.410 4.000 ;
    END
  END ch_out[127]
  PIN ch_out[128]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1860.170 56.000 1860.450 60.000 ;
    END
  END ch_out[128]
  PIN ch_out[129]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 842.890 0.000 843.170 4.000 ;
    END
  END ch_out[129]
  PIN ch_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 65.650 0.000 65.930 4.000 ;
    END
  END ch_out[12]
  PIN ch_out[130]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1865.610 56.000 1865.890 60.000 ;
    END
  END ch_out[130]
  PIN ch_out[131]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 864.650 0.000 864.930 4.000 ;
    END
  END ch_out[131]
  PIN ch_out[132]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1871.050 56.000 1871.330 60.000 ;
    END
  END ch_out[132]
  PIN ch_out[133]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 886.410 0.000 886.690 4.000 ;
    END
  END ch_out[133]
  PIN ch_out[134]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1876.490 56.000 1876.770 60.000 ;
    END
  END ch_out[134]
  PIN ch_out[135]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 908.170 0.000 908.450 4.000 ;
    END
  END ch_out[135]
  PIN ch_out[136]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1881.930 56.000 1882.210 60.000 ;
    END
  END ch_out[136]
  PIN ch_out[137]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 929.930 0.000 930.210 4.000 ;
    END
  END ch_out[137]
  PIN ch_out[138]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1887.370 56.000 1887.650 60.000 ;
    END
  END ch_out[138]
  PIN ch_out[139]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 951.690 0.000 951.970 4.000 ;
    END
  END ch_out[139]
  PIN ch_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1035.670 56.000 1035.950 60.000 ;
    END
  END ch_out[13]
  PIN ch_out[140]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1892.810 56.000 1893.090 60.000 ;
    END
  END ch_out[140]
  PIN ch_out[141]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 973.450 0.000 973.730 4.000 ;
    END
  END ch_out[141]
  PIN ch_out[142]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1100.270 0.000 1100.550 4.000 ;
    END
  END ch_out[142]
  PIN ch_out[143]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1111.150 0.000 1111.430 4.000 ;
    END
  END ch_out[143]
  PIN ch_out[144]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1122.030 0.000 1122.310 4.000 ;
    END
  END ch_out[144]
  PIN ch_out[145]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1132.910 0.000 1133.190 4.000 ;
    END
  END ch_out[145]
  PIN ch_out[146]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1143.790 0.000 1144.070 4.000 ;
    END
  END ch_out[146]
  PIN ch_out[147]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1154.670 0.000 1154.950 4.000 ;
    END
  END ch_out[147]
  PIN ch_out[148]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1165.550 0.000 1165.830 4.000 ;
    END
  END ch_out[148]
  PIN ch_out[149]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1176.430 0.000 1176.710 4.000 ;
    END
  END ch_out[149]
  PIN ch_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1038.390 56.000 1038.670 60.000 ;
    END
  END ch_out[14]
  PIN ch_out[150]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1187.310 0.000 1187.590 4.000 ;
    END
  END ch_out[150]
  PIN ch_out[151]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1198.190 0.000 1198.470 4.000 ;
    END
  END ch_out[151]
  PIN ch_out[152]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1209.070 0.000 1209.350 4.000 ;
    END
  END ch_out[152]
  PIN ch_out[153]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1219.950 0.000 1220.230 4.000 ;
    END
  END ch_out[153]
  PIN ch_out[154]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1230.830 0.000 1231.110 4.000 ;
    END
  END ch_out[154]
  PIN ch_out[155]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1241.710 0.000 1241.990 4.000 ;
    END
  END ch_out[155]
  PIN ch_out[156]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1252.590 0.000 1252.870 4.000 ;
    END
  END ch_out[156]
  PIN ch_out[157]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1263.470 0.000 1263.750 4.000 ;
    END
  END ch_out[157]
  PIN ch_out[158]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1274.350 0.000 1274.630 4.000 ;
    END
  END ch_out[158]
  PIN ch_out[159]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1285.230 0.000 1285.510 4.000 ;
    END
  END ch_out[159]
  PIN ch_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1041.110 56.000 1041.390 60.000 ;
    END
  END ch_out[15]
  PIN ch_out[160]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1296.110 0.000 1296.390 4.000 ;
    END
  END ch_out[160]
  PIN ch_out[161]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1306.990 0.000 1307.270 4.000 ;
    END
  END ch_out[161]
  PIN ch_out[162]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1317.870 0.000 1318.150 4.000 ;
    END
  END ch_out[162]
  PIN ch_out[163]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1328.750 0.000 1329.030 4.000 ;
    END
  END ch_out[163]
  PIN ch_out[164]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1339.630 0.000 1339.910 4.000 ;
    END
  END ch_out[164]
  PIN ch_out[165]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1350.510 0.000 1350.790 4.000 ;
    END
  END ch_out[165]
  PIN ch_out[166]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1361.390 0.000 1361.670 4.000 ;
    END
  END ch_out[166]
  PIN ch_out[167]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1372.270 0.000 1372.550 4.000 ;
    END
  END ch_out[167]
  PIN ch_out[168]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1383.150 0.000 1383.430 4.000 ;
    END
  END ch_out[168]
  PIN ch_out[169]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1394.030 0.000 1394.310 4.000 ;
    END
  END ch_out[169]
  PIN ch_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 87.410 0.000 87.690 4.000 ;
    END
  END ch_out[16]
  PIN ch_out[170]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1404.910 0.000 1405.190 4.000 ;
    END
  END ch_out[170]
  PIN ch_out[171]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1415.790 0.000 1416.070 4.000 ;
    END
  END ch_out[171]
  PIN ch_out[172]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1426.670 0.000 1426.950 4.000 ;
    END
  END ch_out[172]
  PIN ch_out[173]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1437.550 0.000 1437.830 4.000 ;
    END
  END ch_out[173]
  PIN ch_out[174]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1448.430 0.000 1448.710 4.000 ;
    END
  END ch_out[174]
  PIN ch_out[175]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1459.310 0.000 1459.590 4.000 ;
    END
  END ch_out[175]
  PIN ch_out[176]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1470.190 0.000 1470.470 4.000 ;
    END
  END ch_out[176]
  PIN ch_out[177]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1481.070 0.000 1481.350 4.000 ;
    END
  END ch_out[177]
  PIN ch_out[178]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1491.950 0.000 1492.230 4.000 ;
    END
  END ch_out[178]
  PIN ch_out[179]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1502.830 0.000 1503.110 4.000 ;
    END
  END ch_out[179]
  PIN ch_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1046.550 56.000 1046.830 60.000 ;
    END
  END ch_out[17]
  PIN ch_out[180]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1513.710 0.000 1513.990 4.000 ;
    END
  END ch_out[180]
  PIN ch_out[181]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1524.590 0.000 1524.870 4.000 ;
    END
  END ch_out[181]
  PIN ch_out[182]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1535.470 0.000 1535.750 4.000 ;
    END
  END ch_out[182]
  PIN ch_out[183]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1546.350 0.000 1546.630 4.000 ;
    END
  END ch_out[183]
  PIN ch_out[184]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1557.230 0.000 1557.510 4.000 ;
    END
  END ch_out[184]
  PIN ch_out[185]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1568.110 0.000 1568.390 4.000 ;
    END
  END ch_out[185]
  PIN ch_out[186]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1578.990 0.000 1579.270 4.000 ;
    END
  END ch_out[186]
  PIN ch_out[187]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1589.870 0.000 1590.150 4.000 ;
    END
  END ch_out[187]
  PIN ch_out[188]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1800.330 0.000 1800.610 4.000 ;
    END
  END ch_out[188]
  PIN ch_out[189]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1811.210 0.000 1811.490 4.000 ;
    END
  END ch_out[189]
  PIN ch_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1049.270 56.000 1049.550 60.000 ;
    END
  END ch_out[18]
  PIN ch_out[190]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1822.090 0.000 1822.370 4.000 ;
    END
  END ch_out[190]
  PIN ch_out[191]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1832.970 0.000 1833.250 4.000 ;
    END
  END ch_out[191]
  PIN ch_out[192]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1843.850 0.000 1844.130 4.000 ;
    END
  END ch_out[192]
  PIN ch_out[193]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1854.730 0.000 1855.010 4.000 ;
    END
  END ch_out[193]
  PIN ch_out[194]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1865.610 0.000 1865.890 4.000 ;
    END
  END ch_out[194]
  PIN ch_out[195]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1876.490 0.000 1876.770 4.000 ;
    END
  END ch_out[195]
  PIN ch_out[196]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1887.370 0.000 1887.650 4.000 ;
    END
  END ch_out[196]
  PIN ch_out[197]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1898.250 0.000 1898.530 4.000 ;
    END
  END ch_out[197]
  PIN ch_out[198]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1909.130 0.000 1909.410 4.000 ;
    END
  END ch_out[198]
  PIN ch_out[199]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1920.010 0.000 1920.290 4.000 ;
    END
  END ch_out[199]
  PIN ch_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1051.990 56.000 1052.270 60.000 ;
    END
  END ch_out[19]
  PIN ch_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1003.030 56.000 1003.310 60.000 ;
    END
  END ch_out[1]
  PIN ch_out[200]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1930.890 0.000 1931.170 4.000 ;
    END
  END ch_out[200]
  PIN ch_out[201]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1941.770 0.000 1942.050 4.000 ;
    END
  END ch_out[201]
  PIN ch_out[202]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1952.650 0.000 1952.930 4.000 ;
    END
  END ch_out[202]
  PIN ch_out[203]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1963.530 0.000 1963.810 4.000 ;
    END
  END ch_out[203]
  PIN ch_out[204]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1974.410 0.000 1974.690 4.000 ;
    END
  END ch_out[204]
  PIN ch_out[205]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1985.290 0.000 1985.570 4.000 ;
    END
  END ch_out[205]
  PIN ch_out[206]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1996.170 0.000 1996.450 4.000 ;
    END
  END ch_out[206]
  PIN ch_out[207]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2007.050 0.000 2007.330 4.000 ;
    END
  END ch_out[207]
  PIN ch_out[208]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2017.930 0.000 2018.210 4.000 ;
    END
  END ch_out[208]
  PIN ch_out[209]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2028.810 0.000 2029.090 4.000 ;
    END
  END ch_out[209]
  PIN ch_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 109.170 0.000 109.450 4.000 ;
    END
  END ch_out[20]
  PIN ch_out[210]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2039.690 0.000 2039.970 4.000 ;
    END
  END ch_out[210]
  PIN ch_out[211]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2050.570 0.000 2050.850 4.000 ;
    END
  END ch_out[211]
  PIN ch_out[212]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2061.450 0.000 2061.730 4.000 ;
    END
  END ch_out[212]
  PIN ch_out[213]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2072.330 0.000 2072.610 4.000 ;
    END
  END ch_out[213]
  PIN ch_out[214]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2083.210 0.000 2083.490 4.000 ;
    END
  END ch_out[214]
  PIN ch_out[215]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2094.090 0.000 2094.370 4.000 ;
    END
  END ch_out[215]
  PIN ch_out[216]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2104.970 0.000 2105.250 4.000 ;
    END
  END ch_out[216]
  PIN ch_out[217]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2115.850 0.000 2116.130 4.000 ;
    END
  END ch_out[217]
  PIN ch_out[218]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2126.730 0.000 2127.010 4.000 ;
    END
  END ch_out[218]
  PIN ch_out[219]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2137.610 0.000 2137.890 4.000 ;
    END
  END ch_out[219]
  PIN ch_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1057.430 56.000 1057.710 60.000 ;
    END
  END ch_out[21]
  PIN ch_out[220]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2148.490 0.000 2148.770 4.000 ;
    END
  END ch_out[220]
  PIN ch_out[221]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2159.370 0.000 2159.650 4.000 ;
    END
  END ch_out[221]
  PIN ch_out[222]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2170.250 0.000 2170.530 4.000 ;
    END
  END ch_out[222]
  PIN ch_out[223]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2181.130 0.000 2181.410 4.000 ;
    END
  END ch_out[223]
  PIN ch_out[224]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2192.010 0.000 2192.290 4.000 ;
    END
  END ch_out[224]
  PIN ch_out[225]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2202.890 0.000 2203.170 4.000 ;
    END
  END ch_out[225]
  PIN ch_out[226]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2213.770 0.000 2214.050 4.000 ;
    END
  END ch_out[226]
  PIN ch_out[227]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2224.650 0.000 2224.930 4.000 ;
    END
  END ch_out[227]
  PIN ch_out[228]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2235.530 0.000 2235.810 4.000 ;
    END
  END ch_out[228]
  PIN ch_out[229]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2246.410 0.000 2246.690 4.000 ;
    END
  END ch_out[229]
  PIN ch_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1060.150 56.000 1060.430 60.000 ;
    END
  END ch_out[22]
  PIN ch_out[230]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2257.290 0.000 2257.570 4.000 ;
    END
  END ch_out[230]
  PIN ch_out[231]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2268.170 0.000 2268.450 4.000 ;
    END
  END ch_out[231]
  PIN ch_out[232]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2279.050 0.000 2279.330 4.000 ;
    END
  END ch_out[232]
  PIN ch_out[233]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2289.930 0.000 2290.210 4.000 ;
    END
  END ch_out[233]
  PIN ch_out[234]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2300.810 0.000 2301.090 4.000 ;
    END
  END ch_out[234]
  PIN ch_out[235]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2311.690 0.000 2311.970 4.000 ;
    END
  END ch_out[235]
  PIN ch_out[236]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2322.570 0.000 2322.850 4.000 ;
    END
  END ch_out[236]
  PIN ch_out[237]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2333.450 0.000 2333.730 4.000 ;
    END
  END ch_out[237]
  PIN ch_out[238]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2344.330 0.000 2344.610 4.000 ;
    END
  END ch_out[238]
  PIN ch_out[239]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2355.210 0.000 2355.490 4.000 ;
    END
  END ch_out[239]
  PIN ch_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1062.870 56.000 1063.150 60.000 ;
    END
  END ch_out[23]
  PIN ch_out[240]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2366.090 0.000 2366.370 4.000 ;
    END
  END ch_out[240]
  PIN ch_out[241]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2376.970 0.000 2377.250 4.000 ;
    END
  END ch_out[241]
  PIN ch_out[242]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2387.850 0.000 2388.130 4.000 ;
    END
  END ch_out[242]
  PIN ch_out[243]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2398.730 0.000 2399.010 4.000 ;
    END
  END ch_out[243]
  PIN ch_out[244]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2409.610 0.000 2409.890 4.000 ;
    END
  END ch_out[244]
  PIN ch_out[245]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2420.490 0.000 2420.770 4.000 ;
    END
  END ch_out[245]
  PIN ch_out[246]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2431.370 0.000 2431.650 4.000 ;
    END
  END ch_out[246]
  PIN ch_out[247]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2442.250 0.000 2442.530 4.000 ;
    END
  END ch_out[247]
  PIN ch_out[248]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2453.130 0.000 2453.410 4.000 ;
    END
  END ch_out[248]
  PIN ch_out[249]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2464.010 0.000 2464.290 4.000 ;
    END
  END ch_out[249]
  PIN ch_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 130.930 0.000 131.210 4.000 ;
    END
  END ch_out[24]
  PIN ch_out[250]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2474.890 0.000 2475.170 4.000 ;
    END
  END ch_out[250]
  PIN ch_out[251]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2485.770 0.000 2486.050 4.000 ;
    END
  END ch_out[251]
  PIN ch_out[252]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 2443.610 56.000 2443.890 60.000 ;
    END
  END ch_out[252]
  PIN ch_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1068.310 56.000 1068.590 60.000 ;
    END
  END ch_out[25]
  PIN ch_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1071.030 56.000 1071.310 60.000 ;
    END
  END ch_out[26]
  PIN ch_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 147.250 0.000 147.530 4.000 ;
    END
  END ch_out[27]
  PIN ch_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1076.470 56.000 1076.750 60.000 ;
    END
  END ch_out[28]
  PIN ch_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1079.190 56.000 1079.470 60.000 ;
    END
  END ch_out[29]
  PIN ch_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 11.250 0.000 11.530 4.000 ;
    END
  END ch_out[2]
  PIN ch_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 163.570 0.000 163.850 4.000 ;
    END
  END ch_out[30]
  PIN ch_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1084.630 56.000 1084.910 60.000 ;
    END
  END ch_out[31]
  PIN ch_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1087.350 56.000 1087.630 60.000 ;
    END
  END ch_out[32]
  PIN ch_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 179.890 0.000 180.170 4.000 ;
    END
  END ch_out[33]
  PIN ch_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1092.790 56.000 1093.070 60.000 ;
    END
  END ch_out[34]
  PIN ch_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1095.510 56.000 1095.790 60.000 ;
    END
  END ch_out[35]
  PIN ch_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 196.210 0.000 196.490 4.000 ;
    END
  END ch_out[36]
  PIN ch_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1100.950 56.000 1101.230 60.000 ;
    END
  END ch_out[37]
  PIN ch_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1103.670 56.000 1103.950 60.000 ;
    END
  END ch_out[38]
  PIN ch_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 212.530 0.000 212.810 4.000 ;
    END
  END ch_out[39]
  PIN ch_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1008.470 56.000 1008.750 60.000 ;
    END
  END ch_out[3]
  PIN ch_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1109.110 56.000 1109.390 60.000 ;
    END
  END ch_out[40]
  PIN ch_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1111.830 56.000 1112.110 60.000 ;
    END
  END ch_out[41]
  PIN ch_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 228.850 0.000 229.130 4.000 ;
    END
  END ch_out[42]
  PIN ch_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1117.270 56.000 1117.550 60.000 ;
    END
  END ch_out[43]
  PIN ch_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1119.990 56.000 1120.270 60.000 ;
    END
  END ch_out[44]
  PIN ch_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 245.170 0.000 245.450 4.000 ;
    END
  END ch_out[45]
  PIN ch_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1125.430 56.000 1125.710 60.000 ;
    END
  END ch_out[46]
  PIN ch_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1128.150 56.000 1128.430 60.000 ;
    END
  END ch_out[47]
  PIN ch_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 261.490 0.000 261.770 4.000 ;
    END
  END ch_out[48]
  PIN ch_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1133.590 56.000 1133.870 60.000 ;
    END
  END ch_out[49]
  PIN ch_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1011.190 56.000 1011.470 60.000 ;
    END
  END ch_out[4]
  PIN ch_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1136.310 56.000 1136.590 60.000 ;
    END
  END ch_out[50]
  PIN ch_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 277.810 0.000 278.090 4.000 ;
    END
  END ch_out[51]
  PIN ch_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1141.750 56.000 1142.030 60.000 ;
    END
  END ch_out[52]
  PIN ch_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1144.470 56.000 1144.750 60.000 ;
    END
  END ch_out[53]
  PIN ch_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 294.130 0.000 294.410 4.000 ;
    END
  END ch_out[54]
  PIN ch_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1149.910 56.000 1150.190 60.000 ;
    END
  END ch_out[55]
  PIN ch_out[56]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1152.630 56.000 1152.910 60.000 ;
    END
  END ch_out[56]
  PIN ch_out[57]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 310.450 0.000 310.730 4.000 ;
    END
  END ch_out[57]
  PIN ch_out[58]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1158.070 56.000 1158.350 60.000 ;
    END
  END ch_out[58]
  PIN ch_out[59]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1160.790 56.000 1161.070 60.000 ;
    END
  END ch_out[59]
  PIN ch_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1013.910 56.000 1014.190 60.000 ;
    END
  END ch_out[5]
  PIN ch_out[60]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 326.770 0.000 327.050 4.000 ;
    END
  END ch_out[60]
  PIN ch_out[61]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1166.230 56.000 1166.510 60.000 ;
    END
  END ch_out[61]
  PIN ch_out[62]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1168.950 56.000 1169.230 60.000 ;
    END
  END ch_out[62]
  PIN ch_out[63]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 343.090 0.000 343.370 4.000 ;
    END
  END ch_out[63]
  PIN ch_out[64]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1174.390 56.000 1174.670 60.000 ;
    END
  END ch_out[64]
  PIN ch_out[65]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1177.110 56.000 1177.390 60.000 ;
    END
  END ch_out[65]
  PIN ch_out[66]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 359.410 0.000 359.690 4.000 ;
    END
  END ch_out[66]
  PIN ch_out[67]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1182.550 56.000 1182.830 60.000 ;
    END
  END ch_out[67]
  PIN ch_out[68]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1185.270 56.000 1185.550 60.000 ;
    END
  END ch_out[68]
  PIN ch_out[69]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 375.730 0.000 376.010 4.000 ;
    END
  END ch_out[69]
  PIN ch_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1016.630 56.000 1016.910 60.000 ;
    END
  END ch_out[6]
  PIN ch_out[70]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1190.710 56.000 1190.990 60.000 ;
    END
  END ch_out[70]
  PIN ch_out[71]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1193.430 56.000 1193.710 60.000 ;
    END
  END ch_out[71]
  PIN ch_out[72]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 392.050 0.000 392.330 4.000 ;
    END
  END ch_out[72]
  PIN ch_out[73]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1198.870 56.000 1199.150 60.000 ;
    END
  END ch_out[73]
  PIN ch_out[74]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1201.590 56.000 1201.870 60.000 ;
    END
  END ch_out[74]
  PIN ch_out[75]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 408.370 0.000 408.650 4.000 ;
    END
  END ch_out[75]
  PIN ch_out[76]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1207.030 56.000 1207.310 60.000 ;
    END
  END ch_out[76]
  PIN ch_out[77]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1209.750 56.000 1210.030 60.000 ;
    END
  END ch_out[77]
  PIN ch_out[78]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 424.690 0.000 424.970 4.000 ;
    END
  END ch_out[78]
  PIN ch_out[79]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1215.190 56.000 1215.470 60.000 ;
    END
  END ch_out[79]
  PIN ch_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1019.350 56.000 1019.630 60.000 ;
    END
  END ch_out[7]
  PIN ch_out[80]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1217.910 56.000 1218.190 60.000 ;
    END
  END ch_out[80]
  PIN ch_out[81]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 441.010 0.000 441.290 4.000 ;
    END
  END ch_out[81]
  PIN ch_out[82]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1223.350 56.000 1223.630 60.000 ;
    END
  END ch_out[82]
  PIN ch_out[83]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1226.070 56.000 1226.350 60.000 ;
    END
  END ch_out[83]
  PIN ch_out[84]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END ch_out[84]
  PIN ch_out[85]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1231.510 56.000 1231.790 60.000 ;
    END
  END ch_out[85]
  PIN ch_out[86]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1234.230 56.000 1234.510 60.000 ;
    END
  END ch_out[86]
  PIN ch_out[87]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 473.650 0.000 473.930 4.000 ;
    END
  END ch_out[87]
  PIN ch_out[88]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1239.670 56.000 1239.950 60.000 ;
    END
  END ch_out[88]
  PIN ch_out[89]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1242.390 56.000 1242.670 60.000 ;
    END
  END ch_out[89]
  PIN ch_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 43.890 0.000 44.170 4.000 ;
    END
  END ch_out[8]
  PIN ch_out[90]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 489.970 0.000 490.250 4.000 ;
    END
  END ch_out[90]
  PIN ch_out[91]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1247.830 56.000 1248.110 60.000 ;
    END
  END ch_out[91]
  PIN ch_out[92]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1250.550 56.000 1250.830 60.000 ;
    END
  END ch_out[92]
  PIN ch_out[93]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 506.290 0.000 506.570 4.000 ;
    END
  END ch_out[93]
  PIN ch_out[94]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1255.990 56.000 1256.270 60.000 ;
    END
  END ch_out[94]
  PIN ch_out[95]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1258.710 56.000 1258.990 60.000 ;
    END
  END ch_out[95]
  PIN ch_out[96]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 522.610 0.000 522.890 4.000 ;
    END
  END ch_out[96]
  PIN ch_out[97]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1264.150 56.000 1264.430 60.000 ;
    END
  END ch_out[97]
  PIN ch_out[98]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1266.870 56.000 1267.150 60.000 ;
    END
  END ch_out[98]
  PIN ch_out[99]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 538.930 0.000 539.210 4.000 ;
    END
  END ch_out[99]
  PIN ch_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 1024.790 56.000 1025.070 60.000 ;
    END
  END ch_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met2 ;
        RECT -2.080 3.280 -0.480 56.560 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.080 3.280 2651.680 4.880 ;
    END
    PORT
      LAYER met3 ;
        RECT -2.080 54.960 2651.680 56.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 2650.080 3.280 2651.680 56.560 ;
    END
    PORT
      LAYER met2 ;
        RECT 334.540 -0.020 336.140 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 994.180 -0.020 995.780 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1653.820 -0.020 1655.420 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 2313.460 -0.020 2315.060 59.860 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 14.840 2654.980 16.440 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 24.360 2654.980 25.960 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 33.880 2654.980 35.480 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 43.400 2654.980 45.000 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT -5.380 -0.020 -3.780 59.860 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 -0.020 2654.980 1.580 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 58.260 2654.980 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 2653.380 -0.020 2654.980 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 337.840 -0.020 339.440 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 997.480 -0.020 999.080 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 1657.120 -0.020 1658.720 59.860 ;
    END
    PORT
      LAYER met2 ;
        RECT 2316.760 -0.020 2318.360 59.860 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 18.140 2654.980 19.740 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 27.660 2654.980 29.260 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 37.180 2654.980 38.780 ;
    END
    PORT
      LAYER met3 ;
        RECT -5.380 46.700 2654.980 48.300 ;
    END
  END vssd1
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 2644.080 49.045 ;
      LAYER met1 ;
        RECT 0.650 55.720 1000.030 59.800 ;
        RECT 1000.870 55.720 1002.750 59.800 ;
        RECT 1003.590 55.720 1005.470 59.800 ;
        RECT 1006.310 55.720 1008.190 59.800 ;
        RECT 1009.030 55.720 1010.910 59.800 ;
        RECT 1011.750 55.720 1013.630 59.800 ;
        RECT 1014.470 55.720 1016.350 59.800 ;
        RECT 1017.190 55.720 1019.070 59.800 ;
        RECT 1019.910 55.720 1021.790 59.800 ;
        RECT 1022.630 55.720 1024.510 59.800 ;
        RECT 1025.350 55.720 1027.230 59.800 ;
        RECT 1028.070 55.720 1029.950 59.800 ;
        RECT 1030.790 55.720 1032.670 59.800 ;
        RECT 1033.510 55.720 1035.390 59.800 ;
        RECT 1036.230 55.720 1038.110 59.800 ;
        RECT 1038.950 55.720 1040.830 59.800 ;
        RECT 1041.670 55.720 1043.550 59.800 ;
        RECT 1044.390 55.720 1046.270 59.800 ;
        RECT 1047.110 55.720 1048.990 59.800 ;
        RECT 1049.830 55.720 1051.710 59.800 ;
        RECT 1052.550 55.720 1054.430 59.800 ;
        RECT 1055.270 55.720 1057.150 59.800 ;
        RECT 1057.990 55.720 1059.870 59.800 ;
        RECT 1060.710 55.720 1062.590 59.800 ;
        RECT 1063.430 55.720 1065.310 59.800 ;
        RECT 1066.150 55.720 1068.030 59.800 ;
        RECT 1068.870 55.720 1070.750 59.800 ;
        RECT 1071.590 55.720 1073.470 59.800 ;
        RECT 1074.310 55.720 1076.190 59.800 ;
        RECT 1077.030 55.720 1078.910 59.800 ;
        RECT 1079.750 55.720 1081.630 59.800 ;
        RECT 1082.470 55.720 1084.350 59.800 ;
        RECT 1085.190 55.720 1087.070 59.800 ;
        RECT 1087.910 55.720 1089.790 59.800 ;
        RECT 1090.630 55.720 1092.510 59.800 ;
        RECT 1093.350 55.720 1095.230 59.800 ;
        RECT 1096.070 55.720 1097.950 59.800 ;
        RECT 1098.790 55.720 1100.670 59.800 ;
        RECT 1101.510 55.720 1103.390 59.800 ;
        RECT 1104.230 55.720 1106.110 59.800 ;
        RECT 1106.950 55.720 1108.830 59.800 ;
        RECT 1109.670 55.720 1111.550 59.800 ;
        RECT 1112.390 55.720 1114.270 59.800 ;
        RECT 1115.110 55.720 1116.990 59.800 ;
        RECT 1117.830 55.720 1119.710 59.800 ;
        RECT 1120.550 55.720 1122.430 59.800 ;
        RECT 1123.270 55.720 1125.150 59.800 ;
        RECT 1125.990 55.720 1127.870 59.800 ;
        RECT 1128.710 55.720 1130.590 59.800 ;
        RECT 1131.430 55.720 1133.310 59.800 ;
        RECT 1134.150 55.720 1136.030 59.800 ;
        RECT 1136.870 55.720 1138.750 59.800 ;
        RECT 1139.590 55.720 1141.470 59.800 ;
        RECT 1142.310 55.720 1144.190 59.800 ;
        RECT 1145.030 55.720 1146.910 59.800 ;
        RECT 1147.750 55.720 1149.630 59.800 ;
        RECT 1150.470 55.720 1152.350 59.800 ;
        RECT 1153.190 55.720 1155.070 59.800 ;
        RECT 1155.910 55.720 1157.790 59.800 ;
        RECT 1158.630 55.720 1160.510 59.800 ;
        RECT 1161.350 55.720 1163.230 59.800 ;
        RECT 1164.070 55.720 1165.950 59.800 ;
        RECT 1166.790 55.720 1168.670 59.800 ;
        RECT 1169.510 55.720 1171.390 59.800 ;
        RECT 1172.230 55.720 1174.110 59.800 ;
        RECT 1174.950 55.720 1176.830 59.800 ;
        RECT 1177.670 55.720 1179.550 59.800 ;
        RECT 1180.390 55.720 1182.270 59.800 ;
        RECT 1183.110 55.720 1184.990 59.800 ;
        RECT 1185.830 55.720 1187.710 59.800 ;
        RECT 1188.550 55.720 1190.430 59.800 ;
        RECT 1191.270 55.720 1193.150 59.800 ;
        RECT 1193.990 55.720 1195.870 59.800 ;
        RECT 1196.710 55.720 1198.590 59.800 ;
        RECT 1199.430 55.720 1201.310 59.800 ;
        RECT 1202.150 55.720 1204.030 59.800 ;
        RECT 1204.870 55.720 1206.750 59.800 ;
        RECT 1207.590 55.720 1209.470 59.800 ;
        RECT 1210.310 55.720 1212.190 59.800 ;
        RECT 1213.030 55.720 1214.910 59.800 ;
        RECT 1215.750 55.720 1217.630 59.800 ;
        RECT 1218.470 55.720 1220.350 59.800 ;
        RECT 0.650 55.580 1220.350 55.720 ;
        RECT 1221.190 55.720 1223.070 59.800 ;
        RECT 1223.910 55.720 1225.790 59.800 ;
        RECT 1226.630 55.720 1228.510 59.800 ;
        RECT 1229.350 55.720 1231.230 59.800 ;
        RECT 1232.070 55.720 1233.950 59.800 ;
        RECT 1234.790 55.720 1236.670 59.800 ;
        RECT 1237.510 55.720 1239.390 59.800 ;
        RECT 1240.230 55.720 1242.110 59.800 ;
        RECT 1242.950 55.720 1244.830 59.800 ;
        RECT 1245.670 55.720 1247.550 59.800 ;
        RECT 1248.390 55.720 1250.270 59.800 ;
        RECT 1251.110 55.720 1252.990 59.800 ;
        RECT 1253.830 55.720 1255.710 59.800 ;
        RECT 1256.550 55.720 1258.430 59.800 ;
        RECT 1259.270 55.720 1261.150 59.800 ;
        RECT 1261.990 55.720 1263.870 59.800 ;
        RECT 1264.710 55.720 1266.590 59.800 ;
        RECT 1267.430 55.720 1269.310 59.800 ;
        RECT 1270.150 55.720 1272.030 59.800 ;
        RECT 1272.870 55.720 1274.750 59.800 ;
        RECT 1275.590 55.720 1277.470 59.800 ;
        RECT 1278.310 55.720 1280.190 59.800 ;
        RECT 1281.030 55.720 1282.910 59.800 ;
        RECT 1283.750 55.720 1285.630 59.800 ;
        RECT 1286.470 55.720 1800.050 59.800 ;
        RECT 1800.890 55.720 1802.770 59.800 ;
        RECT 1803.610 55.720 1805.490 59.800 ;
        RECT 1806.330 55.720 1808.210 59.800 ;
        RECT 1809.050 55.720 1810.930 59.800 ;
        RECT 1811.770 55.720 1813.650 59.800 ;
        RECT 1814.490 55.720 1816.370 59.800 ;
        RECT 1817.210 55.720 1819.090 59.800 ;
        RECT 1819.930 55.720 1821.810 59.800 ;
        RECT 1822.650 55.720 1824.530 59.800 ;
        RECT 1825.370 55.720 1827.250 59.800 ;
        RECT 1828.090 55.720 1829.970 59.800 ;
        RECT 1830.810 55.720 1832.690 59.800 ;
        RECT 1833.530 55.720 1835.410 59.800 ;
        RECT 1836.250 55.720 1838.130 59.800 ;
        RECT 1838.970 55.720 1840.850 59.800 ;
        RECT 1841.690 55.720 1843.570 59.800 ;
        RECT 1844.410 55.720 1846.290 59.800 ;
        RECT 1847.130 55.720 1849.010 59.800 ;
        RECT 1849.850 55.720 1851.730 59.800 ;
        RECT 1852.570 55.720 1854.450 59.800 ;
        RECT 1855.290 55.720 1857.170 59.800 ;
        RECT 1858.010 55.720 1859.890 59.800 ;
        RECT 1860.730 55.720 1862.610 59.800 ;
        RECT 1863.450 55.720 1865.330 59.800 ;
        RECT 1866.170 55.720 1868.050 59.800 ;
        RECT 1868.890 55.720 1870.770 59.800 ;
        RECT 1871.610 55.720 1873.490 59.800 ;
        RECT 1874.330 55.720 1876.210 59.800 ;
        RECT 1877.050 55.720 1878.930 59.800 ;
        RECT 1879.770 55.720 1881.650 59.800 ;
        RECT 1882.490 55.720 1884.370 59.800 ;
        RECT 1885.210 55.720 1887.090 59.800 ;
        RECT 1887.930 55.720 1889.810 59.800 ;
        RECT 1890.650 55.720 1892.530 59.800 ;
        RECT 1893.370 55.720 1895.250 59.800 ;
        RECT 1896.090 55.720 1897.970 59.800 ;
        RECT 1898.810 55.720 1900.690 59.800 ;
        RECT 1901.530 55.720 1903.410 59.800 ;
        RECT 1904.250 55.720 1906.130 59.800 ;
        RECT 1906.970 55.720 1908.850 59.800 ;
        RECT 1909.690 55.720 1911.570 59.800 ;
        RECT 1912.410 55.720 1914.290 59.800 ;
        RECT 1915.130 55.720 1917.010 59.800 ;
        RECT 1917.850 55.720 1919.730 59.800 ;
        RECT 1920.570 55.720 1922.450 59.800 ;
        RECT 1221.190 55.580 1922.450 55.720 ;
        RECT 1923.290 55.720 1925.170 59.800 ;
        RECT 1926.010 55.720 1927.890 59.800 ;
        RECT 1928.730 55.720 1930.610 59.800 ;
        RECT 1931.450 55.720 1933.330 59.800 ;
        RECT 1934.170 55.720 1936.050 59.800 ;
        RECT 1936.890 55.720 1938.770 59.800 ;
        RECT 1939.610 55.720 1941.490 59.800 ;
        RECT 1942.330 55.720 1944.210 59.800 ;
        RECT 1945.050 55.720 1946.930 59.800 ;
        RECT 1947.770 55.720 1949.650 59.800 ;
        RECT 1950.490 55.720 1952.370 59.800 ;
        RECT 1953.210 55.720 1955.090 59.800 ;
        RECT 1955.930 55.720 1957.810 59.800 ;
        RECT 1958.650 55.720 1960.530 59.800 ;
        RECT 1961.370 55.720 1963.250 59.800 ;
        RECT 1964.090 55.720 1965.970 59.800 ;
        RECT 1966.810 55.720 1968.690 59.800 ;
        RECT 1969.530 55.720 1971.410 59.800 ;
        RECT 1972.250 55.720 1974.130 59.800 ;
        RECT 1974.970 55.720 1976.850 59.800 ;
        RECT 1977.690 55.720 1979.570 59.800 ;
        RECT 1980.410 55.720 1982.290 59.800 ;
        RECT 1983.130 55.720 1985.010 59.800 ;
        RECT 1923.290 55.580 1985.010 55.720 ;
        RECT 1985.850 55.720 1987.730 59.800 ;
        RECT 1988.570 55.720 1990.450 59.800 ;
        RECT 1991.290 55.720 1993.170 59.800 ;
        RECT 1994.010 55.720 1995.890 59.800 ;
        RECT 1996.730 55.720 1998.610 59.800 ;
        RECT 1999.450 55.720 2001.330 59.800 ;
        RECT 2002.170 55.720 2004.050 59.800 ;
        RECT 2004.890 55.720 2006.770 59.800 ;
        RECT 2007.610 55.720 2009.490 59.800 ;
        RECT 2010.330 55.720 2012.210 59.800 ;
        RECT 2013.050 55.720 2014.930 59.800 ;
        RECT 2015.770 55.720 2017.650 59.800 ;
        RECT 2018.490 55.720 2020.370 59.800 ;
        RECT 2021.210 55.720 2199.890 59.800 ;
        RECT 2200.730 55.720 2201.250 59.800 ;
        RECT 2202.090 55.720 2202.610 59.800 ;
        RECT 2203.450 55.720 2203.970 59.800 ;
        RECT 2204.810 55.720 2205.330 59.800 ;
        RECT 2206.170 55.720 2206.690 59.800 ;
        RECT 2207.530 55.720 2208.050 59.800 ;
        RECT 2208.890 55.720 2209.410 59.800 ;
        RECT 2210.250 55.720 2210.770 59.800 ;
        RECT 2211.610 55.720 2212.130 59.800 ;
        RECT 2212.970 55.720 2213.490 59.800 ;
        RECT 1985.850 55.580 2213.490 55.720 ;
        RECT 2214.330 55.720 2214.850 59.800 ;
        RECT 2215.690 55.720 2216.210 59.800 ;
        RECT 2217.050 55.720 2217.570 59.800 ;
        RECT 2218.410 55.720 2218.930 59.800 ;
        RECT 2219.770 55.720 2220.290 59.800 ;
        RECT 2221.130 55.720 2221.650 59.800 ;
        RECT 2222.490 55.720 2223.010 59.800 ;
        RECT 2223.850 55.720 2224.370 59.800 ;
        RECT 2225.210 55.720 2225.730 59.800 ;
        RECT 2226.570 55.720 2227.090 59.800 ;
        RECT 2227.930 55.720 2228.450 59.800 ;
        RECT 2229.290 55.720 2229.810 59.800 ;
        RECT 2230.650 55.720 2231.170 59.800 ;
        RECT 2232.010 55.720 2232.530 59.800 ;
        RECT 2233.370 55.720 2233.890 59.800 ;
        RECT 2234.730 55.720 2235.250 59.800 ;
        RECT 2214.330 55.580 2235.250 55.720 ;
        RECT 2236.090 55.720 2236.610 59.800 ;
        RECT 2237.450 55.720 2237.970 59.800 ;
        RECT 2238.810 55.720 2239.330 59.800 ;
        RECT 2240.170 55.720 2240.690 59.800 ;
        RECT 2241.530 55.720 2242.050 59.800 ;
        RECT 2242.890 55.720 2399.810 59.800 ;
        RECT 2400.650 55.720 2401.170 59.800 ;
        RECT 2236.090 55.580 2401.170 55.720 ;
        RECT 2402.010 55.720 2402.530 59.800 ;
        RECT 2403.370 55.720 2403.890 59.800 ;
        RECT 2404.730 55.720 2405.250 59.800 ;
        RECT 2406.090 55.720 2406.610 59.800 ;
        RECT 2407.450 55.720 2407.970 59.800 ;
        RECT 2408.810 55.720 2409.330 59.800 ;
        RECT 2410.170 55.720 2410.690 59.800 ;
        RECT 2411.530 55.720 2412.050 59.800 ;
        RECT 2412.890 55.720 2413.410 59.800 ;
        RECT 2414.250 55.720 2414.770 59.800 ;
        RECT 2402.010 55.580 2414.770 55.720 ;
        RECT 2415.610 55.720 2416.130 59.800 ;
        RECT 2416.970 55.720 2417.490 59.800 ;
        RECT 2418.330 55.720 2418.850 59.800 ;
        RECT 2419.690 55.720 2420.210 59.800 ;
        RECT 2421.050 55.720 2421.570 59.800 ;
        RECT 2422.410 55.720 2422.930 59.800 ;
        RECT 2423.770 55.720 2424.290 59.800 ;
        RECT 2425.130 55.720 2425.650 59.800 ;
        RECT 2426.490 55.720 2427.010 59.800 ;
        RECT 2427.850 55.720 2428.370 59.800 ;
        RECT 2429.210 55.720 2429.730 59.800 ;
        RECT 2430.570 55.720 2431.090 59.800 ;
        RECT 2431.930 55.720 2432.450 59.800 ;
        RECT 2433.290 55.720 2433.810 59.800 ;
        RECT 2434.650 55.720 2435.170 59.800 ;
        RECT 2436.010 55.720 2436.530 59.800 ;
        RECT 2437.370 55.720 2437.890 59.800 ;
        RECT 2438.730 55.720 2439.250 59.800 ;
        RECT 2440.090 55.720 2440.610 59.800 ;
        RECT 2441.450 55.720 2441.970 59.800 ;
        RECT 2442.810 55.720 2443.330 59.800 ;
        RECT 2444.170 55.720 2644.080 59.800 ;
        RECT 2415.610 55.580 2644.080 55.720 ;
        RECT 0.650 4.280 2644.080 55.580 ;
        RECT 0.930 0.040 5.530 4.280 ;
        RECT 6.370 0.040 10.970 4.280 ;
        RECT 11.810 0.040 16.410 4.280 ;
        RECT 17.250 0.040 21.850 4.280 ;
        RECT 22.690 0.040 27.290 4.280 ;
        RECT 28.130 0.040 32.730 4.280 ;
        RECT 33.570 0.040 38.170 4.280 ;
        RECT 39.010 0.040 43.610 4.280 ;
        RECT 44.450 0.040 49.050 4.280 ;
        RECT 49.890 0.040 54.490 4.280 ;
        RECT 55.330 0.040 59.930 4.280 ;
        RECT 60.770 0.040 65.370 4.280 ;
        RECT 66.210 0.040 70.810 4.280 ;
        RECT 71.650 0.040 76.250 4.280 ;
        RECT 77.090 0.040 81.690 4.280 ;
        RECT 82.530 0.040 87.130 4.280 ;
        RECT 87.970 0.040 92.570 4.280 ;
        RECT 93.410 0.040 98.010 4.280 ;
        RECT 98.850 0.040 103.450 4.280 ;
        RECT 104.290 0.040 108.890 4.280 ;
        RECT 109.730 0.040 114.330 4.280 ;
        RECT 115.170 0.040 119.770 4.280 ;
        RECT 120.610 0.040 125.210 4.280 ;
        RECT 126.050 0.040 130.650 4.280 ;
        RECT 131.490 0.040 136.090 4.280 ;
        RECT 136.930 0.040 141.530 4.280 ;
        RECT 142.370 0.040 146.970 4.280 ;
        RECT 147.810 0.040 152.410 4.280 ;
        RECT 153.250 0.040 157.850 4.280 ;
        RECT 158.690 0.040 163.290 4.280 ;
        RECT 164.130 0.040 168.730 4.280 ;
        RECT 169.570 0.040 174.170 4.280 ;
        RECT 175.010 0.040 179.610 4.280 ;
        RECT 180.450 0.040 185.050 4.280 ;
        RECT 185.890 0.040 190.490 4.280 ;
        RECT 191.330 0.040 195.930 4.280 ;
        RECT 196.770 0.040 201.370 4.280 ;
        RECT 202.210 0.040 206.810 4.280 ;
        RECT 207.650 0.040 212.250 4.280 ;
        RECT 213.090 0.040 217.690 4.280 ;
        RECT 218.530 0.040 223.130 4.280 ;
        RECT 223.970 0.040 228.570 4.280 ;
        RECT 229.410 0.040 234.010 4.280 ;
        RECT 234.850 0.040 239.450 4.280 ;
        RECT 240.290 0.040 244.890 4.280 ;
        RECT 245.730 0.040 250.330 4.280 ;
        RECT 251.170 0.040 255.770 4.280 ;
        RECT 256.610 0.040 261.210 4.280 ;
        RECT 262.050 0.040 266.650 4.280 ;
        RECT 267.490 0.040 272.090 4.280 ;
        RECT 272.930 0.040 277.530 4.280 ;
        RECT 278.370 0.040 282.970 4.280 ;
        RECT 283.810 0.040 288.410 4.280 ;
        RECT 289.250 0.040 293.850 4.280 ;
        RECT 294.690 0.040 299.290 4.280 ;
        RECT 300.130 0.040 304.730 4.280 ;
        RECT 305.570 0.040 310.170 4.280 ;
        RECT 311.010 0.040 315.610 4.280 ;
        RECT 316.450 0.040 321.050 4.280 ;
        RECT 321.890 0.040 326.490 4.280 ;
        RECT 327.330 0.040 331.930 4.280 ;
        RECT 332.770 0.040 337.370 4.280 ;
        RECT 338.210 0.040 342.810 4.280 ;
        RECT 343.650 0.040 348.250 4.280 ;
        RECT 349.090 0.040 353.690 4.280 ;
        RECT 354.530 0.040 359.130 4.280 ;
        RECT 359.970 0.040 364.570 4.280 ;
        RECT 365.410 0.040 370.010 4.280 ;
        RECT 370.850 0.040 375.450 4.280 ;
        RECT 376.290 0.040 380.890 4.280 ;
        RECT 381.730 0.040 386.330 4.280 ;
        RECT 387.170 0.040 391.770 4.280 ;
        RECT 392.610 0.040 397.210 4.280 ;
        RECT 398.050 0.040 402.650 4.280 ;
        RECT 403.490 0.040 408.090 4.280 ;
        RECT 408.930 0.040 413.530 4.280 ;
        RECT 414.370 0.040 418.970 4.280 ;
        RECT 419.810 0.040 424.410 4.280 ;
        RECT 425.250 0.040 429.850 4.280 ;
        RECT 430.690 0.040 435.290 4.280 ;
        RECT 436.130 0.040 440.730 4.280 ;
        RECT 441.570 0.040 446.170 4.280 ;
        RECT 447.010 0.040 451.610 4.280 ;
        RECT 452.450 0.040 457.050 4.280 ;
        RECT 457.890 0.040 462.490 4.280 ;
        RECT 463.330 0.040 467.930 4.280 ;
        RECT 468.770 0.040 473.370 4.280 ;
        RECT 474.210 0.040 478.810 4.280 ;
        RECT 479.650 0.040 484.250 4.280 ;
        RECT 485.090 0.040 489.690 4.280 ;
        RECT 490.530 0.040 495.130 4.280 ;
        RECT 495.970 0.040 500.570 4.280 ;
        RECT 501.410 0.040 506.010 4.280 ;
        RECT 506.850 0.040 511.450 4.280 ;
        RECT 512.290 0.040 516.890 4.280 ;
        RECT 517.730 0.040 522.330 4.280 ;
        RECT 523.170 0.040 527.770 4.280 ;
        RECT 528.610 0.040 533.210 4.280 ;
        RECT 534.050 0.040 538.650 4.280 ;
        RECT 539.490 0.040 544.090 4.280 ;
        RECT 544.930 0.040 549.530 4.280 ;
        RECT 550.370 0.040 554.970 4.280 ;
        RECT 555.810 0.040 560.410 4.280 ;
        RECT 561.250 0.040 565.850 4.280 ;
        RECT 566.690 0.040 571.290 4.280 ;
        RECT 572.130 0.040 599.850 4.280 ;
        RECT 600.690 0.040 610.730 4.280 ;
        RECT 611.570 0.040 621.610 4.280 ;
        RECT 622.450 0.040 632.490 4.280 ;
        RECT 633.330 0.040 643.370 4.280 ;
        RECT 644.210 0.040 654.250 4.280 ;
        RECT 655.090 0.040 665.130 4.280 ;
        RECT 665.970 0.040 676.010 4.280 ;
        RECT 676.850 0.040 686.890 4.280 ;
        RECT 687.730 0.040 697.770 4.280 ;
        RECT 698.610 0.040 708.650 4.280 ;
        RECT 709.490 0.040 719.530 4.280 ;
        RECT 720.370 0.040 730.410 4.280 ;
        RECT 731.250 0.040 741.290 4.280 ;
        RECT 742.130 0.040 752.170 4.280 ;
        RECT 753.010 0.040 763.050 4.280 ;
        RECT 763.890 0.040 773.930 4.280 ;
        RECT 774.770 0.040 784.810 4.280 ;
        RECT 785.650 0.040 795.690 4.280 ;
        RECT 796.530 0.040 806.570 4.280 ;
        RECT 807.410 0.040 809.970 4.280 ;
        RECT 810.810 0.040 820.850 4.280 ;
        RECT 821.690 0.040 831.730 4.280 ;
        RECT 832.570 0.040 842.610 4.280 ;
        RECT 843.450 0.040 853.490 4.280 ;
        RECT 854.330 0.040 864.370 4.280 ;
        RECT 865.210 0.040 875.250 4.280 ;
        RECT 876.090 0.040 886.130 4.280 ;
        RECT 886.970 0.040 897.010 4.280 ;
        RECT 897.850 0.040 907.890 4.280 ;
        RECT 908.730 0.040 918.770 4.280 ;
        RECT 919.610 0.040 929.650 4.280 ;
        RECT 930.490 0.040 940.530 4.280 ;
        RECT 941.370 0.040 951.410 4.280 ;
        RECT 952.250 0.040 962.290 4.280 ;
        RECT 963.130 0.040 973.170 4.280 ;
        RECT 974.010 0.040 1099.990 4.280 ;
        RECT 1100.830 0.040 1110.870 4.280 ;
        RECT 1111.710 0.040 1121.750 4.280 ;
        RECT 1122.590 0.040 1132.630 4.280 ;
        RECT 1133.470 0.040 1143.510 4.280 ;
        RECT 1144.350 0.040 1154.390 4.280 ;
        RECT 1155.230 0.040 1165.270 4.280 ;
        RECT 1166.110 0.040 1176.150 4.280 ;
        RECT 1176.990 0.040 1187.030 4.280 ;
        RECT 1187.870 0.040 1197.910 4.280 ;
        RECT 1198.750 0.040 1208.790 4.280 ;
        RECT 1209.630 0.040 1219.670 4.280 ;
        RECT 1220.510 0.040 1230.550 4.280 ;
        RECT 1231.390 0.040 1241.430 4.280 ;
        RECT 1242.270 0.040 1252.310 4.280 ;
        RECT 1253.150 0.040 1263.190 4.280 ;
        RECT 1264.030 0.040 1274.070 4.280 ;
        RECT 1274.910 0.040 1284.950 4.280 ;
        RECT 1285.790 0.040 1295.830 4.280 ;
        RECT 1296.670 0.040 1306.710 4.280 ;
        RECT 1307.550 0.040 1317.590 4.280 ;
        RECT 1318.430 0.040 1328.470 4.280 ;
        RECT 1329.310 0.040 1339.350 4.280 ;
        RECT 1340.190 0.040 1350.230 4.280 ;
        RECT 1351.070 0.040 1361.110 4.280 ;
        RECT 1361.950 0.040 1371.990 4.280 ;
        RECT 1372.830 0.040 1382.870 4.280 ;
        RECT 1383.710 0.040 1393.750 4.280 ;
        RECT 1394.590 0.040 1404.630 4.280 ;
        RECT 1405.470 0.040 1415.510 4.280 ;
        RECT 1416.350 0.040 1426.390 4.280 ;
        RECT 1427.230 0.040 1437.270 4.280 ;
        RECT 1438.110 0.040 1448.150 4.280 ;
        RECT 1448.990 0.040 1459.030 4.280 ;
        RECT 1459.870 0.040 1469.910 4.280 ;
        RECT 1470.750 0.040 1480.790 4.280 ;
        RECT 1481.630 0.040 1491.670 4.280 ;
        RECT 1492.510 0.040 1502.550 4.280 ;
        RECT 1503.390 0.040 1513.430 4.280 ;
        RECT 1514.270 0.040 1524.310 4.280 ;
        RECT 1525.150 0.040 1535.190 4.280 ;
        RECT 1536.030 0.040 1546.070 4.280 ;
        RECT 1546.910 0.040 1556.950 4.280 ;
        RECT 1557.790 0.040 1567.830 4.280 ;
        RECT 1568.670 0.040 1578.710 4.280 ;
        RECT 1579.550 0.040 1589.590 4.280 ;
        RECT 1590.430 0.040 1800.050 4.280 ;
        RECT 1800.890 0.040 1810.930 4.280 ;
        RECT 1811.770 0.040 1821.810 4.280 ;
        RECT 1822.650 0.040 1832.690 4.280 ;
        RECT 1833.530 0.040 1843.570 4.280 ;
        RECT 1844.410 0.040 1854.450 4.280 ;
        RECT 1855.290 0.040 1865.330 4.280 ;
        RECT 1866.170 0.040 1876.210 4.280 ;
        RECT 1877.050 0.040 1887.090 4.280 ;
        RECT 1887.930 0.040 1897.970 4.280 ;
        RECT 1898.810 0.040 1908.850 4.280 ;
        RECT 1909.690 0.040 1919.730 4.280 ;
        RECT 1920.570 0.040 1930.610 4.280 ;
        RECT 1931.450 0.040 1941.490 4.280 ;
        RECT 1942.330 0.040 1952.370 4.280 ;
        RECT 1953.210 0.040 1963.250 4.280 ;
        RECT 1964.090 0.040 1974.130 4.280 ;
        RECT 1974.970 0.040 1985.010 4.280 ;
        RECT 1985.850 0.040 1995.890 4.280 ;
        RECT 1996.730 0.040 2006.770 4.280 ;
        RECT 2007.610 0.040 2017.650 4.280 ;
        RECT 2018.490 0.040 2028.530 4.280 ;
        RECT 2029.370 0.040 2039.410 4.280 ;
        RECT 2040.250 0.040 2050.290 4.280 ;
        RECT 2051.130 0.040 2061.170 4.280 ;
        RECT 2062.010 0.040 2072.050 4.280 ;
        RECT 2072.890 0.040 2082.930 4.280 ;
        RECT 2083.770 0.040 2093.810 4.280 ;
        RECT 2094.650 0.040 2104.690 4.280 ;
        RECT 2105.530 0.040 2115.570 4.280 ;
        RECT 2116.410 0.040 2126.450 4.280 ;
        RECT 2127.290 0.040 2137.330 4.280 ;
        RECT 2138.170 0.040 2148.210 4.280 ;
        RECT 2149.050 0.040 2159.090 4.280 ;
        RECT 2159.930 0.040 2169.970 4.280 ;
        RECT 2170.810 0.040 2180.850 4.280 ;
        RECT 2181.690 0.040 2191.730 4.280 ;
        RECT 2192.570 0.040 2202.610 4.280 ;
        RECT 2203.450 0.040 2213.490 4.280 ;
        RECT 2214.330 0.040 2224.370 4.280 ;
        RECT 2225.210 0.040 2235.250 4.280 ;
        RECT 2236.090 0.040 2246.130 4.280 ;
        RECT 2246.970 0.040 2257.010 4.280 ;
        RECT 2257.850 0.040 2267.890 4.280 ;
        RECT 2268.730 0.040 2278.770 4.280 ;
        RECT 2279.610 0.040 2289.650 4.280 ;
        RECT 2290.490 0.040 2300.530 4.280 ;
        RECT 2301.370 0.040 2311.410 4.280 ;
        RECT 2312.250 0.040 2322.290 4.280 ;
        RECT 2323.130 0.040 2333.170 4.280 ;
        RECT 2334.010 0.040 2344.050 4.280 ;
        RECT 2344.890 0.040 2354.930 4.280 ;
        RECT 2355.770 0.040 2365.810 4.280 ;
        RECT 2366.650 0.040 2376.690 4.280 ;
        RECT 2377.530 0.040 2387.570 4.280 ;
        RECT 2388.410 0.040 2398.450 4.280 ;
        RECT 2399.290 0.040 2409.330 4.280 ;
        RECT 2410.170 0.040 2420.210 4.280 ;
        RECT 2421.050 0.040 2431.090 4.280 ;
        RECT 2431.930 0.040 2441.970 4.280 ;
        RECT 2442.810 0.040 2452.850 4.280 ;
        RECT 2453.690 0.040 2463.730 4.280 ;
        RECT 2464.570 0.040 2474.610 4.280 ;
        RECT 2475.450 0.040 2485.490 4.280 ;
        RECT 2486.330 0.040 2496.370 4.280 ;
        RECT 2497.210 0.040 2644.080 4.280 ;
      LAYER met2 ;
        RECT 4.240 0.010 334.260 59.830 ;
        RECT 336.420 0.010 337.560 59.830 ;
        RECT 339.720 0.010 993.900 59.830 ;
        RECT 996.060 0.010 997.200 59.830 ;
        RECT 999.360 0.010 1653.540 59.830 ;
        RECT 1655.700 0.010 1656.840 59.830 ;
        RECT 1659.000 0.010 2313.180 59.830 ;
        RECT 2315.340 0.010 2316.480 59.830 ;
        RECT 2318.640 0.010 2571.300 59.830 ;
      LAYER met3 ;
        RECT 141.745 56.960 1970.115 57.625 ;
        RECT 141.745 48.700 1970.115 54.560 ;
        RECT 141.745 45.400 1970.115 46.300 ;
        RECT 141.745 39.180 1970.115 43.000 ;
        RECT 141.745 35.880 1970.115 36.780 ;
        RECT 141.745 29.660 1970.115 33.480 ;
        RECT 141.745 26.360 1970.115 27.260 ;
        RECT 141.745 20.140 1970.115 23.960 ;
        RECT 141.745 16.840 1970.115 17.740 ;
        RECT 141.745 5.280 1970.115 14.440 ;
        RECT 141.745 2.215 1970.115 2.880 ;
  END
END bus_rep_south
END LIBRARY

