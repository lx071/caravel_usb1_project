// This is the unpowered netlist.
module pinmux_top (cfg_dco_mode,
    cfg_pll_enb,
    cfg_strap_pad_ctrl,
    cpu_clk,
    cpu_intf_rst_n,
    e_reset_n,
    i2cm_clk_i,
    i2cm_clk_o,
    i2cm_clk_oen,
    i2cm_data_i,
    i2cm_data_o,
    i2cm_data_oen,
    i2cm_intr,
    i2cm_rst_n,
    int_pll_clock,
    ir_intr,
    ir_rx,
    ir_tx,
    mclk,
    p_reset_n,
    pll_ref_clk,
    pulse1m_mclk,
    qspim_rst_n,
    reg_ack,
    reg_cs,
    reg_peri_ack,
    reg_peri_cs,
    reg_peri_wr,
    reg_wr,
    riscv_tck,
    riscv_tdi,
    riscv_tdo,
    riscv_tdo_en,
    riscv_tms,
    riscv_trst_n,
    rtc_clk,
    rtc_intr,
    s_reset_n,
    sflash_sck,
    sm_a1,
    sm_a2,
    sm_b1,
    sm_b2,
    soft_irq,
    spim_miso,
    spim_mosi,
    spim_sck,
    spis_miso,
    spis_mosi,
    spis_sck,
    spis_ssn,
    sspim_rst_n,
    uartm_rxd,
    uartm_txd,
    usb_clk,
    usb_dn_i,
    usb_dn_o,
    usb_dp_i,
    usb_dp_o,
    usb_intr,
    usb_oen,
    usb_rst_n,
    user_clock1,
    user_clock2,
    wbd_clk_int,
    wbd_clk_pinmux,
    xtal_clk,
    cfg_cska_pinmux,
    cfg_dc_trim,
    cfg_pll_fed_div,
    cfg_riscv_ctrl,
    cpu_core_rst_n,
    digital_io_in,
    digital_io_oen,
    digital_io_out,
    irq_lines,
    pinmux_debug,
    reg_addr,
    reg_be,
    reg_peri_addr,
    reg_peri_be,
    reg_peri_rdata,
    reg_peri_wdata,
    reg_rdata,
    reg_wdata,
    sflash_di,
    sflash_do,
    sflash_oen,
    sflash_ss,
    spim_ssn,
    strap_sticky,
    strap_uartm,
    system_strap,
    uart_rst_n,
    uart_rxd,
    uart_txd,
    user_irq);
 output cfg_dco_mode;
 output cfg_pll_enb;
 input cfg_strap_pad_ctrl;
 input cpu_clk;
 output cpu_intf_rst_n;
 input e_reset_n;
 output i2cm_clk_i;
 input i2cm_clk_o;
 input i2cm_clk_oen;
 output i2cm_data_i;
 input i2cm_data_o;
 input i2cm_data_oen;
 input i2cm_intr;
 output i2cm_rst_n;
 input int_pll_clock;
 input ir_intr;
 output ir_rx;
 input ir_tx;
 input mclk;
 input p_reset_n;
 output pll_ref_clk;
 output pulse1m_mclk;
 output qspim_rst_n;
 output reg_ack;
 input reg_cs;
 input reg_peri_ack;
 output reg_peri_cs;
 output reg_peri_wr;
 input reg_wr;
 output riscv_tck;
 output riscv_tdi;
 input riscv_tdo;
 input riscv_tdo_en;
 output riscv_tms;
 output riscv_trst_n;
 output rtc_clk;
 input rtc_intr;
 input s_reset_n;
 input sflash_sck;
 input sm_a1;
 input sm_a2;
 input sm_b1;
 input sm_b2;
 output soft_irq;
 input spim_miso;
 output spim_mosi;
 input spim_sck;
 input spis_miso;
 output spis_mosi;
 output spis_sck;
 output spis_ssn;
 output sspim_rst_n;
 output uartm_rxd;
 input uartm_txd;
 output usb_clk;
 output usb_dn_i;
 input usb_dn_o;
 output usb_dp_i;
 input usb_dp_o;
 input usb_intr;
 input usb_oen;
 output usb_rst_n;
 input user_clock1;
 input user_clock2;
 input wbd_clk_int;
 output wbd_clk_pinmux;
 output xtal_clk;
 input [3:0] cfg_cska_pinmux;
 output [25:0] cfg_dc_trim;
 output [4:0] cfg_pll_fed_div;
 output [15:0] cfg_riscv_ctrl;
 output [3:0] cpu_core_rst_n;
 input [37:0] digital_io_in;
 output [37:0] digital_io_oen;
 output [37:0] digital_io_out;
 output [31:0] irq_lines;
 output [31:0] pinmux_debug;
 input [10:0] reg_addr;
 input [3:0] reg_be;
 output [10:0] reg_peri_addr;
 output [3:0] reg_peri_be;
 input [31:0] reg_peri_rdata;
 output [31:0] reg_peri_wdata;
 output [31:0] reg_rdata;
 input [31:0] reg_wdata;
 output [3:0] sflash_di;
 input [3:0] sflash_do;
 input [3:0] sflash_oen;
 input [3:0] sflash_ss;
 input [3:0] spim_ssn;
 output [31:0] strap_sticky;
 output [1:0] strap_uartm;
 input [31:0] system_strap;
 output [1:0] uart_rst_n;
 output [1:0] uart_rxd;
 input [1:0] uart_txd;
 output [2:0] user_irq;

 wire net1657;
 wire net1667;
 wire net1668;
 wire net1669;
 wire net1670;
 wire net1671;
 wire net1672;
 wire net1673;
 wire net1674;
 wire net1675;
 wire net1676;
 wire net1658;
 wire net1677;
 wire net1678;
 wire net1679;
 wire net1680;
 wire net1681;
 wire net1682;
 wire net1683;
 wire net1684;
 wire net1685;
 wire net1686;
 wire net1659;
 wire net1687;
 wire net1688;
 wire net1660;
 wire net1661;
 wire net1662;
 wire net1663;
 wire net1664;
 wire net1665;
 wire net1666;
 wire _00000_;
 wire _00001_;
 wire _00002_;
 wire _00003_;
 wire _00004_;
 wire _00005_;
 wire _00006_;
 wire _00007_;
 wire _00008_;
 wire _00009_;
 wire _00010_;
 wire _00011_;
 wire _00012_;
 wire _00013_;
 wire _00014_;
 wire _00015_;
 wire _00016_;
 wire _00017_;
 wire _00018_;
 wire _00019_;
 wire _00020_;
 wire _00021_;
 wire _00022_;
 wire _00023_;
 wire _00024_;
 wire _00025_;
 wire _00026_;
 wire _00027_;
 wire _00028_;
 wire _00029_;
 wire _00030_;
 wire _00031_;
 wire _00032_;
 wire _00033_;
 wire _00034_;
 wire _00035_;
 wire _00036_;
 wire _00037_;
 wire _00038_;
 wire _00039_;
 wire _00040_;
 wire _00041_;
 wire _00042_;
 wire _00043_;
 wire _00044_;
 wire _00045_;
 wire _00046_;
 wire _00047_;
 wire _00048_;
 wire _00049_;
 wire _00050_;
 wire _00051_;
 wire _00052_;
 wire _00053_;
 wire _00054_;
 wire _00055_;
 wire _00056_;
 wire _00057_;
 wire _00058_;
 wire _00059_;
 wire _00060_;
 wire _00061_;
 wire _00062_;
 wire _00063_;
 wire _00064_;
 wire _00065_;
 wire _00066_;
 wire _00067_;
 wire _00068_;
 wire _00069_;
 wire _00070_;
 wire _00071_;
 wire _00072_;
 wire _00073_;
 wire _00074_;
 wire _00075_;
 wire _00076_;
 wire _00077_;
 wire _00078_;
 wire _00079_;
 wire _00080_;
 wire _00081_;
 wire _00082_;
 wire _00083_;
 wire _00084_;
 wire _00085_;
 wire _00086_;
 wire _00087_;
 wire _00088_;
 wire _00089_;
 wire _00090_;
 wire _00091_;
 wire _00092_;
 wire _00093_;
 wire _00094_;
 wire _00095_;
 wire _00096_;
 wire _00097_;
 wire _00098_;
 wire _00099_;
 wire _00100_;
 wire _00101_;
 wire _00102_;
 wire _00103_;
 wire _00104_;
 wire _00105_;
 wire _00106_;
 wire _00107_;
 wire _00108_;
 wire _00109_;
 wire _00110_;
 wire _00111_;
 wire _00112_;
 wire _00113_;
 wire _00114_;
 wire _00115_;
 wire _00116_;
 wire _00117_;
 wire _00118_;
 wire _00119_;
 wire _00120_;
 wire _00121_;
 wire _00122_;
 wire _00123_;
 wire _00124_;
 wire _00125_;
 wire _00126_;
 wire _00127_;
 wire _00128_;
 wire _00129_;
 wire _00130_;
 wire _00131_;
 wire _00132_;
 wire _00133_;
 wire _00134_;
 wire _00135_;
 wire _00136_;
 wire _00137_;
 wire _00138_;
 wire _00139_;
 wire _00140_;
 wire _00141_;
 wire _00142_;
 wire _00143_;
 wire _00144_;
 wire _00145_;
 wire _00146_;
 wire _00147_;
 wire _00148_;
 wire _00149_;
 wire _00150_;
 wire _00151_;
 wire _00152_;
 wire _00153_;
 wire _00154_;
 wire _00155_;
 wire _00156_;
 wire _00157_;
 wire _00158_;
 wire _00159_;
 wire _00160_;
 wire _00161_;
 wire _00162_;
 wire _00163_;
 wire _00164_;
 wire _00165_;
 wire _00166_;
 wire _00167_;
 wire _00168_;
 wire _00169_;
 wire _00170_;
 wire _00171_;
 wire _00172_;
 wire _00173_;
 wire _00174_;
 wire _00175_;
 wire _00176_;
 wire _00177_;
 wire _00178_;
 wire _00179_;
 wire _00180_;
 wire _00181_;
 wire _00182_;
 wire _00183_;
 wire _00184_;
 wire _00185_;
 wire _00186_;
 wire _00187_;
 wire _00188_;
 wire _00189_;
 wire _00190_;
 wire _00191_;
 wire _00192_;
 wire _00193_;
 wire _00194_;
 wire _00195_;
 wire _00196_;
 wire _00197_;
 wire _00198_;
 wire _00199_;
 wire _00200_;
 wire _00201_;
 wire _00202_;
 wire _00203_;
 wire _00204_;
 wire _00205_;
 wire _00206_;
 wire _00207_;
 wire _00208_;
 wire _00209_;
 wire _00210_;
 wire _00211_;
 wire _00212_;
 wire _00213_;
 wire _00214_;
 wire _00215_;
 wire _00216_;
 wire _00217_;
 wire _00218_;
 wire _00219_;
 wire _00220_;
 wire _00221_;
 wire _00222_;
 wire _00223_;
 wire _00224_;
 wire _00225_;
 wire _00226_;
 wire _00227_;
 wire _00228_;
 wire _00229_;
 wire _00230_;
 wire _00231_;
 wire _00232_;
 wire _00233_;
 wire _00234_;
 wire _00235_;
 wire _00236_;
 wire _00237_;
 wire _00238_;
 wire _00239_;
 wire _00240_;
 wire _00241_;
 wire _00242_;
 wire _00243_;
 wire _00244_;
 wire _00245_;
 wire _00246_;
 wire _00247_;
 wire _00248_;
 wire _00249_;
 wire _00250_;
 wire _00251_;
 wire _00252_;
 wire _00253_;
 wire _00254_;
 wire _00255_;
 wire _00256_;
 wire _00257_;
 wire _00258_;
 wire _00259_;
 wire _00260_;
 wire _00261_;
 wire _00262_;
 wire _00263_;
 wire _00264_;
 wire _00265_;
 wire _00266_;
 wire _00267_;
 wire _00268_;
 wire _00269_;
 wire _00270_;
 wire _00271_;
 wire _00272_;
 wire _00273_;
 wire _00274_;
 wire _00275_;
 wire _00276_;
 wire _00277_;
 wire _00278_;
 wire _00279_;
 wire _00280_;
 wire _00281_;
 wire _00282_;
 wire _00283_;
 wire _00284_;
 wire _00285_;
 wire _00286_;
 wire _00287_;
 wire _00288_;
 wire _00289_;
 wire _00290_;
 wire _00291_;
 wire _00292_;
 wire _00293_;
 wire _00294_;
 wire _00295_;
 wire _00296_;
 wire _00297_;
 wire _00298_;
 wire _00299_;
 wire _00300_;
 wire _00301_;
 wire _00302_;
 wire _00303_;
 wire _00304_;
 wire _00305_;
 wire _00306_;
 wire _00307_;
 wire _00308_;
 wire _00309_;
 wire _00310_;
 wire _00311_;
 wire _00312_;
 wire _00313_;
 wire _00314_;
 wire _00315_;
 wire _00316_;
 wire _00317_;
 wire _00318_;
 wire _00319_;
 wire _00320_;
 wire _00321_;
 wire _00322_;
 wire _00323_;
 wire _00324_;
 wire _00325_;
 wire _00326_;
 wire _00327_;
 wire _00328_;
 wire _00329_;
 wire _00330_;
 wire _00331_;
 wire _00332_;
 wire _00333_;
 wire _00334_;
 wire _00335_;
 wire _00336_;
 wire _00337_;
 wire _00338_;
 wire _00339_;
 wire _00340_;
 wire _00341_;
 wire _00342_;
 wire _00343_;
 wire _00344_;
 wire _00345_;
 wire _00346_;
 wire _00347_;
 wire _00348_;
 wire _00349_;
 wire _00350_;
 wire _00351_;
 wire _00352_;
 wire _00353_;
 wire _00354_;
 wire _00355_;
 wire _00356_;
 wire _00357_;
 wire _00358_;
 wire _00359_;
 wire _00360_;
 wire _00361_;
 wire _00362_;
 wire _00363_;
 wire _00364_;
 wire _00365_;
 wire _00366_;
 wire _00367_;
 wire _00368_;
 wire _00369_;
 wire _00370_;
 wire _00371_;
 wire _00372_;
 wire _00373_;
 wire _00374_;
 wire _00375_;
 wire _00376_;
 wire _00377_;
 wire _00378_;
 wire _00379_;
 wire _00380_;
 wire _00381_;
 wire _00382_;
 wire _00383_;
 wire _00384_;
 wire _00385_;
 wire _00386_;
 wire _00387_;
 wire _00388_;
 wire _00389_;
 wire _00390_;
 wire _00391_;
 wire _00392_;
 wire _00393_;
 wire _00394_;
 wire _00395_;
 wire _00396_;
 wire _00397_;
 wire _00398_;
 wire _00399_;
 wire _00400_;
 wire _00401_;
 wire _00402_;
 wire _00403_;
 wire _00404_;
 wire _00405_;
 wire _00406_;
 wire _00407_;
 wire _00408_;
 wire _00409_;
 wire _00410_;
 wire _00411_;
 wire _00412_;
 wire _00413_;
 wire _00414_;
 wire _00415_;
 wire _00416_;
 wire _00417_;
 wire _00418_;
 wire _00419_;
 wire _00420_;
 wire _00421_;
 wire _00422_;
 wire _00423_;
 wire _00424_;
 wire _00425_;
 wire _00426_;
 wire _00427_;
 wire _00428_;
 wire _00429_;
 wire _00430_;
 wire _00431_;
 wire _00432_;
 wire _00433_;
 wire _00434_;
 wire _00435_;
 wire _00436_;
 wire _00437_;
 wire _00438_;
 wire _00439_;
 wire _00440_;
 wire _00441_;
 wire _00442_;
 wire _00443_;
 wire _00444_;
 wire _00445_;
 wire _00446_;
 wire _00447_;
 wire _00448_;
 wire _00449_;
 wire _00450_;
 wire _00451_;
 wire _00452_;
 wire _00453_;
 wire _00454_;
 wire _00455_;
 wire _00456_;
 wire _00457_;
 wire _00458_;
 wire _00459_;
 wire _00460_;
 wire _00461_;
 wire _00462_;
 wire _00463_;
 wire _00464_;
 wire _00465_;
 wire _00466_;
 wire _00467_;
 wire _00468_;
 wire _00469_;
 wire _00470_;
 wire _00471_;
 wire _00472_;
 wire _00473_;
 wire _00474_;
 wire _00475_;
 wire _00476_;
 wire _00477_;
 wire _00478_;
 wire _00479_;
 wire _00480_;
 wire _00481_;
 wire _00482_;
 wire _00483_;
 wire _00484_;
 wire _00485_;
 wire _00486_;
 wire _00487_;
 wire _00488_;
 wire _00489_;
 wire _00490_;
 wire _00491_;
 wire _00492_;
 wire _00493_;
 wire _00494_;
 wire _00495_;
 wire _00496_;
 wire _00497_;
 wire _00498_;
 wire _00499_;
 wire _00500_;
 wire _00501_;
 wire _00502_;
 wire _00503_;
 wire _00504_;
 wire _00505_;
 wire _00506_;
 wire _00507_;
 wire _00508_;
 wire _00509_;
 wire _00510_;
 wire _00511_;
 wire _00512_;
 wire _00513_;
 wire _00514_;
 wire _00515_;
 wire _00516_;
 wire _00517_;
 wire _00518_;
 wire _00519_;
 wire _00520_;
 wire _00521_;
 wire _00522_;
 wire _00523_;
 wire _00524_;
 wire _00525_;
 wire _00526_;
 wire _00527_;
 wire _00528_;
 wire _00529_;
 wire _00530_;
 wire _00531_;
 wire _00532_;
 wire _00533_;
 wire _00534_;
 wire _00535_;
 wire _00536_;
 wire _00537_;
 wire _00538_;
 wire _00539_;
 wire _00540_;
 wire _00541_;
 wire _00542_;
 wire _00543_;
 wire _00544_;
 wire _00545_;
 wire _00546_;
 wire _00547_;
 wire _00548_;
 wire _00549_;
 wire _00550_;
 wire _00551_;
 wire _00552_;
 wire _00553_;
 wire _00554_;
 wire _00555_;
 wire _00556_;
 wire _00557_;
 wire _00558_;
 wire _00559_;
 wire _00560_;
 wire _00561_;
 wire _00562_;
 wire _00563_;
 wire _00564_;
 wire _00565_;
 wire _00566_;
 wire _00567_;
 wire _00568_;
 wire _00569_;
 wire _00570_;
 wire _00571_;
 wire _00572_;
 wire _00573_;
 wire _00574_;
 wire _00575_;
 wire _00576_;
 wire _00577_;
 wire _00578_;
 wire _00579_;
 wire _00580_;
 wire _00581_;
 wire _00582_;
 wire _00583_;
 wire _00584_;
 wire _00585_;
 wire _00586_;
 wire _00587_;
 wire _00588_;
 wire _00589_;
 wire _00590_;
 wire _00591_;
 wire _00592_;
 wire _00593_;
 wire _00594_;
 wire _00595_;
 wire _00596_;
 wire _00597_;
 wire _00598_;
 wire _00599_;
 wire _00600_;
 wire _00601_;
 wire _00602_;
 wire _00603_;
 wire _00604_;
 wire _00605_;
 wire _00606_;
 wire _00607_;
 wire _00608_;
 wire _00609_;
 wire _00610_;
 wire _00611_;
 wire _00612_;
 wire _00613_;
 wire _00614_;
 wire _00615_;
 wire _00616_;
 wire _00617_;
 wire _00618_;
 wire _00619_;
 wire _00620_;
 wire _00621_;
 wire _00622_;
 wire _00623_;
 wire _00624_;
 wire _00625_;
 wire _00626_;
 wire _00627_;
 wire _00628_;
 wire _00629_;
 wire _00630_;
 wire _00631_;
 wire _00632_;
 wire _00633_;
 wire _00634_;
 wire _00635_;
 wire _00636_;
 wire _00637_;
 wire _00638_;
 wire _00639_;
 wire _00640_;
 wire _00641_;
 wire _00642_;
 wire _00643_;
 wire _00644_;
 wire _00645_;
 wire _00646_;
 wire _00647_;
 wire _00648_;
 wire _00649_;
 wire _00650_;
 wire _00651_;
 wire _00652_;
 wire _00653_;
 wire _00654_;
 wire _00655_;
 wire _00656_;
 wire _00657_;
 wire _00658_;
 wire _00659_;
 wire _00660_;
 wire _00661_;
 wire _00662_;
 wire _00663_;
 wire _00664_;
 wire _00665_;
 wire _00666_;
 wire _00667_;
 wire _00668_;
 wire _00669_;
 wire _00670_;
 wire _00671_;
 wire _00672_;
 wire _00673_;
 wire _00674_;
 wire _00675_;
 wire _00676_;
 wire _00677_;
 wire _00678_;
 wire _00679_;
 wire _00680_;
 wire _00681_;
 wire _00682_;
 wire _00683_;
 wire _00684_;
 wire _00685_;
 wire _00686_;
 wire _00687_;
 wire _00688_;
 wire _00689_;
 wire _00690_;
 wire _00691_;
 wire _00692_;
 wire _00693_;
 wire _00694_;
 wire _00695_;
 wire _00696_;
 wire _00697_;
 wire _00698_;
 wire _00699_;
 wire _00700_;
 wire _00701_;
 wire _00702_;
 wire _00703_;
 wire _00704_;
 wire _00705_;
 wire _00706_;
 wire _00707_;
 wire _00708_;
 wire _00709_;
 wire _00710_;
 wire _00711_;
 wire _00712_;
 wire _00713_;
 wire _00714_;
 wire _00715_;
 wire _00716_;
 wire _00717_;
 wire _00718_;
 wire _00719_;
 wire _00720_;
 wire _00721_;
 wire _00722_;
 wire _00723_;
 wire _00724_;
 wire _00725_;
 wire _00726_;
 wire _00727_;
 wire _00728_;
 wire _00729_;
 wire _00730_;
 wire _00731_;
 wire _00732_;
 wire _00733_;
 wire _00734_;
 wire _00735_;
 wire _00736_;
 wire _00737_;
 wire _00738_;
 wire _00739_;
 wire _00740_;
 wire _00741_;
 wire _00742_;
 wire _00743_;
 wire _00744_;
 wire _00745_;
 wire _00746_;
 wire _00747_;
 wire _00748_;
 wire _00749_;
 wire _00750_;
 wire _00751_;
 wire _00752_;
 wire _00753_;
 wire _00754_;
 wire _00755_;
 wire _00756_;
 wire _00757_;
 wire _00758_;
 wire _00759_;
 wire _00760_;
 wire _00761_;
 wire _00762_;
 wire _00763_;
 wire _00764_;
 wire _00765_;
 wire _00766_;
 wire _00767_;
 wire _00768_;
 wire _00769_;
 wire _00770_;
 wire _00771_;
 wire _00772_;
 wire _00773_;
 wire _00774_;
 wire _00775_;
 wire _00776_;
 wire _00777_;
 wire _00778_;
 wire _00779_;
 wire _00780_;
 wire _00781_;
 wire _00782_;
 wire _00783_;
 wire _00784_;
 wire _00785_;
 wire _00786_;
 wire _00787_;
 wire _00788_;
 wire _00789_;
 wire _00790_;
 wire _00791_;
 wire _00792_;
 wire _00793_;
 wire _00794_;
 wire _00795_;
 wire _00796_;
 wire _00797_;
 wire _00798_;
 wire _00799_;
 wire _00800_;
 wire _00801_;
 wire _00802_;
 wire _00803_;
 wire _00804_;
 wire _00805_;
 wire _00806_;
 wire _00807_;
 wire _00808_;
 wire _00809_;
 wire _00810_;
 wire _00811_;
 wire _00812_;
 wire _00813_;
 wire _00814_;
 wire _00815_;
 wire _00816_;
 wire _00817_;
 wire _00818_;
 wire _00819_;
 wire _00820_;
 wire _00821_;
 wire _00822_;
 wire _00823_;
 wire _00824_;
 wire _00825_;
 wire _00826_;
 wire _00827_;
 wire _00828_;
 wire _00829_;
 wire _00830_;
 wire _00831_;
 wire _00832_;
 wire _00833_;
 wire _00834_;
 wire _00835_;
 wire _00836_;
 wire _00837_;
 wire _00838_;
 wire _00839_;
 wire _00840_;
 wire _00841_;
 wire _00842_;
 wire _00843_;
 wire _00844_;
 wire _00845_;
 wire _00846_;
 wire _00847_;
 wire _00848_;
 wire _00849_;
 wire _00850_;
 wire _00851_;
 wire _00852_;
 wire _00853_;
 wire _00854_;
 wire _00855_;
 wire _00856_;
 wire _00857_;
 wire _00858_;
 wire _00859_;
 wire _00860_;
 wire _00861_;
 wire _00862_;
 wire _00863_;
 wire _00864_;
 wire _00865_;
 wire _00866_;
 wire _00867_;
 wire _00868_;
 wire _00869_;
 wire _00870_;
 wire _00871_;
 wire _00872_;
 wire _00873_;
 wire _00874_;
 wire _00875_;
 wire _00876_;
 wire _00877_;
 wire _00878_;
 wire _00879_;
 wire _00880_;
 wire _00881_;
 wire _00882_;
 wire _00883_;
 wire _00884_;
 wire _00885_;
 wire _00886_;
 wire _00887_;
 wire _00888_;
 wire _00889_;
 wire _00890_;
 wire _00891_;
 wire _00892_;
 wire _00893_;
 wire _00894_;
 wire _00895_;
 wire _00896_;
 wire _00897_;
 wire _00898_;
 wire _00899_;
 wire _00900_;
 wire _00901_;
 wire _00902_;
 wire _00903_;
 wire _00904_;
 wire _00905_;
 wire _00906_;
 wire _00907_;
 wire _00908_;
 wire _00909_;
 wire _00910_;
 wire _00911_;
 wire _00912_;
 wire _00913_;
 wire _00914_;
 wire _00915_;
 wire _00916_;
 wire _00917_;
 wire _00918_;
 wire _00919_;
 wire _00920_;
 wire _00921_;
 wire _00922_;
 wire _00923_;
 wire _00924_;
 wire _00925_;
 wire _00926_;
 wire _00927_;
 wire _00928_;
 wire _00929_;
 wire _00930_;
 wire _00931_;
 wire _00932_;
 wire _00933_;
 wire _00934_;
 wire _00935_;
 wire _00936_;
 wire _00937_;
 wire _00938_;
 wire _00939_;
 wire _00940_;
 wire _00941_;
 wire _00942_;
 wire _00943_;
 wire _00944_;
 wire _00945_;
 wire _00946_;
 wire _00947_;
 wire _00948_;
 wire _00949_;
 wire _00950_;
 wire _00951_;
 wire _00952_;
 wire _00953_;
 wire _00954_;
 wire _00955_;
 wire _00956_;
 wire _00957_;
 wire _00958_;
 wire _00959_;
 wire _00960_;
 wire _00961_;
 wire _00962_;
 wire _00963_;
 wire _00964_;
 wire _00965_;
 wire _00966_;
 wire _00967_;
 wire _00968_;
 wire _00969_;
 wire _00970_;
 wire _00971_;
 wire _00972_;
 wire _00973_;
 wire _00974_;
 wire _00975_;
 wire _00976_;
 wire _00977_;
 wire _00978_;
 wire _00979_;
 wire _00980_;
 wire _00981_;
 wire _00982_;
 wire _00983_;
 wire _00984_;
 wire _00985_;
 wire _00986_;
 wire _00987_;
 wire _00988_;
 wire _00989_;
 wire _00990_;
 wire _00991_;
 wire _00992_;
 wire _00993_;
 wire _00994_;
 wire _00995_;
 wire _00996_;
 wire _00997_;
 wire _00998_;
 wire _00999_;
 wire _01000_;
 wire _01001_;
 wire _01002_;
 wire _01003_;
 wire _01004_;
 wire _01005_;
 wire _01006_;
 wire _01007_;
 wire _01008_;
 wire _01009_;
 wire _01010_;
 wire _01011_;
 wire _01012_;
 wire _01013_;
 wire _01014_;
 wire _01015_;
 wire _01016_;
 wire _01017_;
 wire _01018_;
 wire _01019_;
 wire _01020_;
 wire _01021_;
 wire _01022_;
 wire _01023_;
 wire _01024_;
 wire _01025_;
 wire _01026_;
 wire _01027_;
 wire _01028_;
 wire _01029_;
 wire _01030_;
 wire _01031_;
 wire _01032_;
 wire _01033_;
 wire _01034_;
 wire _01035_;
 wire _01036_;
 wire _01037_;
 wire _01038_;
 wire _01039_;
 wire _01040_;
 wire _01041_;
 wire _01042_;
 wire _01043_;
 wire _01044_;
 wire _01045_;
 wire _01046_;
 wire _01047_;
 wire _01048_;
 wire _01049_;
 wire _01050_;
 wire _01051_;
 wire _01052_;
 wire _01053_;
 wire _01054_;
 wire _01055_;
 wire _01056_;
 wire _01057_;
 wire _01058_;
 wire _01059_;
 wire _01060_;
 wire _01061_;
 wire _01062_;
 wire _01063_;
 wire _01064_;
 wire _01065_;
 wire _01066_;
 wire _01067_;
 wire _01068_;
 wire _01069_;
 wire _01070_;
 wire _01071_;
 wire _01072_;
 wire _01073_;
 wire _01074_;
 wire _01075_;
 wire _01076_;
 wire _01077_;
 wire _01078_;
 wire _01079_;
 wire _01080_;
 wire _01081_;
 wire _01082_;
 wire _01083_;
 wire _01084_;
 wire _01085_;
 wire _01086_;
 wire _01087_;
 wire _01088_;
 wire _01089_;
 wire _01090_;
 wire _01091_;
 wire _01092_;
 wire _01093_;
 wire _01094_;
 wire _01095_;
 wire _01096_;
 wire _01097_;
 wire _01098_;
 wire _01099_;
 wire _01100_;
 wire _01101_;
 wire _01102_;
 wire _01103_;
 wire _01104_;
 wire _01105_;
 wire _01106_;
 wire _01107_;
 wire _01108_;
 wire _01109_;
 wire _01110_;
 wire _01111_;
 wire _01112_;
 wire _01113_;
 wire _01114_;
 wire _01115_;
 wire _01116_;
 wire _01117_;
 wire _01118_;
 wire _01119_;
 wire _01120_;
 wire _01121_;
 wire _01122_;
 wire _01123_;
 wire _01124_;
 wire _01125_;
 wire _01126_;
 wire _01127_;
 wire _01128_;
 wire _01129_;
 wire _01130_;
 wire _01131_;
 wire _01132_;
 wire _01133_;
 wire _01134_;
 wire _01135_;
 wire _01136_;
 wire _01137_;
 wire _01138_;
 wire _01139_;
 wire _01140_;
 wire _01141_;
 wire _01142_;
 wire _01143_;
 wire _01144_;
 wire _01145_;
 wire _01146_;
 wire _01147_;
 wire _01148_;
 wire _01149_;
 wire _01150_;
 wire _01151_;
 wire _01152_;
 wire _01153_;
 wire _01154_;
 wire _01155_;
 wire _01156_;
 wire _01157_;
 wire _01158_;
 wire _01159_;
 wire _01160_;
 wire _01161_;
 wire _01162_;
 wire _01163_;
 wire _01164_;
 wire _01165_;
 wire _01166_;
 wire _01167_;
 wire _01168_;
 wire _01169_;
 wire _01170_;
 wire _01171_;
 wire _01172_;
 wire _01173_;
 wire _01174_;
 wire _01175_;
 wire _01176_;
 wire _01177_;
 wire _01178_;
 wire _01179_;
 wire _01180_;
 wire _01181_;
 wire _01182_;
 wire _01183_;
 wire _01184_;
 wire _01185_;
 wire _01186_;
 wire _01187_;
 wire _01188_;
 wire _01189_;
 wire _01190_;
 wire _01191_;
 wire _01192_;
 wire _01193_;
 wire _01194_;
 wire _01195_;
 wire _01196_;
 wire _01197_;
 wire _01198_;
 wire _01199_;
 wire _01200_;
 wire _01201_;
 wire _01202_;
 wire _01203_;
 wire _01204_;
 wire _01205_;
 wire _01206_;
 wire _01207_;
 wire _01208_;
 wire _01209_;
 wire _01210_;
 wire _01211_;
 wire _01212_;
 wire _01213_;
 wire _01214_;
 wire _01215_;
 wire _01216_;
 wire _01217_;
 wire _01218_;
 wire _01219_;
 wire _01220_;
 wire _01221_;
 wire _01222_;
 wire _01223_;
 wire _01224_;
 wire _01225_;
 wire _01226_;
 wire _01227_;
 wire _01228_;
 wire _01229_;
 wire _01230_;
 wire _01231_;
 wire _01232_;
 wire _01233_;
 wire _01234_;
 wire _01235_;
 wire _01236_;
 wire _01237_;
 wire _01238_;
 wire _01239_;
 wire _01240_;
 wire _01241_;
 wire _01242_;
 wire _01243_;
 wire _01244_;
 wire _01245_;
 wire _01246_;
 wire _01247_;
 wire _01248_;
 wire _01249_;
 wire _01250_;
 wire _01251_;
 wire _01252_;
 wire _01253_;
 wire _01254_;
 wire _01255_;
 wire _01256_;
 wire _01257_;
 wire _01258_;
 wire _01259_;
 wire _01260_;
 wire _01261_;
 wire _01262_;
 wire _01263_;
 wire _01264_;
 wire _01265_;
 wire _01266_;
 wire _01267_;
 wire _01268_;
 wire _01269_;
 wire _01270_;
 wire _01271_;
 wire _01272_;
 wire _01273_;
 wire _01274_;
 wire _01275_;
 wire _01276_;
 wire _01277_;
 wire _01278_;
 wire _01279_;
 wire _01280_;
 wire _01281_;
 wire _01282_;
 wire _01283_;
 wire _01284_;
 wire _01285_;
 wire _01286_;
 wire _01287_;
 wire _01288_;
 wire _01289_;
 wire _01290_;
 wire _01291_;
 wire _01292_;
 wire _01293_;
 wire _01294_;
 wire _01295_;
 wire _01296_;
 wire _01297_;
 wire _01298_;
 wire _01299_;
 wire _01300_;
 wire _01301_;
 wire _01302_;
 wire _01303_;
 wire _01304_;
 wire _01305_;
 wire _01306_;
 wire _01307_;
 wire _01308_;
 wire _01309_;
 wire _01310_;
 wire _01311_;
 wire _01312_;
 wire _01313_;
 wire _01314_;
 wire _01315_;
 wire _01316_;
 wire _01317_;
 wire _01318_;
 wire _01319_;
 wire _01320_;
 wire _01321_;
 wire _01322_;
 wire _01323_;
 wire _01324_;
 wire _01325_;
 wire _01326_;
 wire _01327_;
 wire _01328_;
 wire _01329_;
 wire _01330_;
 wire _01331_;
 wire _01332_;
 wire _01333_;
 wire _01334_;
 wire _01335_;
 wire _01336_;
 wire _01337_;
 wire _01338_;
 wire _01339_;
 wire _01340_;
 wire _01341_;
 wire _01342_;
 wire _01343_;
 wire _01344_;
 wire _01345_;
 wire _01346_;
 wire _01347_;
 wire _01348_;
 wire _01349_;
 wire _01350_;
 wire _01351_;
 wire _01352_;
 wire _01353_;
 wire _01354_;
 wire _01355_;
 wire _01356_;
 wire _01357_;
 wire _01358_;
 wire _01359_;
 wire _01360_;
 wire _01361_;
 wire _01362_;
 wire _01363_;
 wire _01364_;
 wire _01365_;
 wire _01366_;
 wire _01367_;
 wire _01368_;
 wire _01369_;
 wire _01370_;
 wire _01371_;
 wire _01372_;
 wire _01373_;
 wire _01374_;
 wire _01375_;
 wire _01376_;
 wire _01377_;
 wire _01378_;
 wire _01379_;
 wire _01380_;
 wire _01381_;
 wire _01382_;
 wire _01383_;
 wire _01384_;
 wire _01385_;
 wire _01386_;
 wire _01387_;
 wire _01388_;
 wire _01389_;
 wire _01390_;
 wire _01391_;
 wire _01392_;
 wire _01393_;
 wire _01394_;
 wire _01395_;
 wire _01396_;
 wire _01397_;
 wire _01398_;
 wire _01399_;
 wire _01400_;
 wire _01401_;
 wire _01402_;
 wire _01403_;
 wire _01404_;
 wire _01405_;
 wire _01406_;
 wire _01407_;
 wire _01408_;
 wire _01409_;
 wire _01410_;
 wire _01411_;
 wire _01412_;
 wire _01413_;
 wire _01414_;
 wire _01415_;
 wire _01416_;
 wire _01417_;
 wire _01418_;
 wire _01419_;
 wire _01420_;
 wire _01421_;
 wire _01422_;
 wire _01423_;
 wire _01424_;
 wire _01425_;
 wire _01426_;
 wire _01427_;
 wire _01428_;
 wire _01429_;
 wire _01430_;
 wire _01431_;
 wire _01432_;
 wire _01433_;
 wire _01434_;
 wire _01435_;
 wire _01436_;
 wire _01437_;
 wire _01438_;
 wire _01439_;
 wire _01440_;
 wire _01441_;
 wire _01442_;
 wire _01443_;
 wire _01444_;
 wire _01445_;
 wire _01446_;
 wire _01447_;
 wire _01448_;
 wire _01449_;
 wire _01450_;
 wire _01451_;
 wire _01452_;
 wire _01453_;
 wire _01454_;
 wire _01455_;
 wire _01456_;
 wire _01457_;
 wire _01458_;
 wire _01459_;
 wire _01460_;
 wire _01461_;
 wire _01462_;
 wire _01463_;
 wire _01464_;
 wire _01465_;
 wire _01466_;
 wire _01467_;
 wire _01468_;
 wire _01469_;
 wire _01470_;
 wire _01471_;
 wire _01472_;
 wire _01473_;
 wire _01474_;
 wire _01475_;
 wire _01476_;
 wire _01477_;
 wire _01478_;
 wire _01479_;
 wire _01480_;
 wire _01481_;
 wire _01482_;
 wire _01483_;
 wire _01484_;
 wire _01485_;
 wire _01486_;
 wire _01487_;
 wire _01488_;
 wire _01489_;
 wire _01490_;
 wire _01491_;
 wire _01492_;
 wire _01493_;
 wire _01494_;
 wire _01495_;
 wire _01496_;
 wire _01497_;
 wire _01498_;
 wire _01499_;
 wire _01500_;
 wire _01501_;
 wire _01502_;
 wire _01503_;
 wire _01504_;
 wire _01505_;
 wire _01506_;
 wire _01507_;
 wire _01508_;
 wire _01509_;
 wire _01510_;
 wire _01511_;
 wire _01512_;
 wire _01513_;
 wire _01514_;
 wire _01515_;
 wire _01516_;
 wire _01517_;
 wire _01518_;
 wire _01519_;
 wire _01520_;
 wire _01521_;
 wire _01522_;
 wire _01523_;
 wire _01524_;
 wire _01525_;
 wire _01526_;
 wire _01527_;
 wire _01528_;
 wire _01529_;
 wire _01530_;
 wire _01531_;
 wire _01532_;
 wire _01533_;
 wire _01534_;
 wire _01535_;
 wire _01536_;
 wire _01537_;
 wire _01538_;
 wire _01539_;
 wire _01540_;
 wire _01541_;
 wire _01542_;
 wire _01543_;
 wire _01544_;
 wire _01545_;
 wire _01546_;
 wire _01547_;
 wire _01548_;
 wire _01549_;
 wire _01550_;
 wire _01551_;
 wire _01552_;
 wire _01553_;
 wire _01554_;
 wire _01555_;
 wire _01556_;
 wire _01557_;
 wire _01558_;
 wire _01559_;
 wire _01560_;
 wire _01561_;
 wire _01562_;
 wire _01563_;
 wire _01564_;
 wire _01565_;
 wire _01566_;
 wire _01567_;
 wire _01568_;
 wire _01569_;
 wire _01570_;
 wire _01571_;
 wire _01572_;
 wire _01573_;
 wire _01574_;
 wire _01575_;
 wire _01576_;
 wire _01577_;
 wire _01578_;
 wire _01579_;
 wire _01580_;
 wire _01581_;
 wire _01582_;
 wire _01583_;
 wire _01584_;
 wire _01585_;
 wire _01586_;
 wire _01587_;
 wire _01588_;
 wire _01589_;
 wire _01590_;
 wire _01591_;
 wire _01592_;
 wire _01593_;
 wire _01594_;
 wire _01595_;
 wire _01596_;
 wire _01597_;
 wire _01598_;
 wire _01599_;
 wire _01600_;
 wire _01601_;
 wire _01602_;
 wire _01603_;
 wire _01604_;
 wire _01605_;
 wire _01606_;
 wire _01607_;
 wire _01608_;
 wire _01609_;
 wire _01610_;
 wire _01611_;
 wire _01612_;
 wire _01613_;
 wire _01614_;
 wire _01615_;
 wire _01616_;
 wire _01617_;
 wire _01618_;
 wire _01619_;
 wire _01620_;
 wire _01621_;
 wire _01622_;
 wire _01623_;
 wire _01624_;
 wire _01625_;
 wire _01626_;
 wire _01627_;
 wire _01628_;
 wire _01629_;
 wire _01630_;
 wire _01631_;
 wire _01632_;
 wire _01633_;
 wire _01634_;
 wire _01635_;
 wire _01636_;
 wire _01637_;
 wire _01638_;
 wire _01639_;
 wire _01640_;
 wire _01641_;
 wire _01642_;
 wire _01643_;
 wire _01644_;
 wire _01645_;
 wire _01646_;
 wire _01647_;
 wire _01648_;
 wire _01649_;
 wire _01650_;
 wire _01651_;
 wire _01652_;
 wire _01653_;
 wire _01654_;
 wire _01655_;
 wire _01656_;
 wire _01657_;
 wire _01658_;
 wire _01659_;
 wire _01660_;
 wire _01661_;
 wire _01662_;
 wire _01663_;
 wire _01664_;
 wire _01665_;
 wire _01666_;
 wire _01667_;
 wire _01668_;
 wire _01669_;
 wire _01670_;
 wire _01671_;
 wire _01672_;
 wire _01673_;
 wire _01674_;
 wire _01675_;
 wire _01677_;
 wire _01678_;
 wire _01679_;
 wire _01680_;
 wire _01681_;
 wire _01682_;
 wire _01683_;
 wire _01684_;
 wire _01685_;
 wire _01686_;
 wire _01687_;
 wire _01688_;
 wire _01689_;
 wire _01690_;
 wire _01691_;
 wire _01692_;
 wire _01693_;
 wire _01694_;
 wire _01695_;
 wire _01696_;
 wire _01697_;
 wire _01698_;
 wire _01699_;
 wire _01700_;
 wire _01701_;
 wire _01702_;
 wire _01703_;
 wire _01704_;
 wire _01705_;
 wire _01706_;
 wire _01707_;
 wire _01708_;
 wire _01709_;
 wire _01710_;
 wire _01711_;
 wire _01712_;
 wire _01713_;
 wire _01714_;
 wire _01715_;
 wire _01716_;
 wire _01717_;
 wire _01718_;
 wire _01719_;
 wire _01720_;
 wire _01721_;
 wire _01722_;
 wire _01723_;
 wire _01724_;
 wire _01725_;
 wire _01726_;
 wire _01727_;
 wire _01728_;
 wire _01729_;
 wire _01730_;
 wire _01731_;
 wire _01732_;
 wire _01733_;
 wire _01734_;
 wire _01735_;
 wire _01736_;
 wire _01737_;
 wire _01738_;
 wire _01739_;
 wire _01740_;
 wire _01741_;
 wire _01742_;
 wire _01743_;
 wire _01744_;
 wire _01745_;
 wire _01746_;
 wire _01747_;
 wire _01748_;
 wire _01749_;
 wire _01750_;
 wire _01751_;
 wire _01752_;
 wire _01753_;
 wire _01754_;
 wire _01755_;
 wire _01756_;
 wire _01757_;
 wire _01758_;
 wire _01759_;
 wire _01760_;
 wire _01761_;
 wire _01762_;
 wire _01763_;
 wire _01764_;
 wire _01765_;
 wire _01766_;
 wire _01767_;
 wire _01768_;
 wire _01769_;
 wire _01770_;
 wire _01771_;
 wire _01772_;
 wire _01773_;
 wire _01774_;
 wire _01775_;
 wire _01776_;
 wire _01777_;
 wire _01778_;
 wire _01779_;
 wire _01780_;
 wire _01781_;
 wire _01782_;
 wire _01783_;
 wire _01784_;
 wire _01785_;
 wire _01786_;
 wire _01787_;
 wire _01788_;
 wire _01789_;
 wire _01790_;
 wire _01791_;
 wire _01792_;
 wire _01793_;
 wire _01794_;
 wire _01795_;
 wire _01796_;
 wire _01797_;
 wire _01798_;
 wire _01799_;
 wire _01800_;
 wire _01801_;
 wire _01802_;
 wire _01803_;
 wire _01804_;
 wire _01805_;
 wire _01806_;
 wire _01807_;
 wire _01808_;
 wire _01809_;
 wire _01810_;
 wire _01811_;
 wire _01812_;
 wire _01813_;
 wire _01814_;
 wire _01815_;
 wire _01816_;
 wire _01817_;
 wire _01818_;
 wire _01819_;
 wire _01820_;
 wire _01821_;
 wire _01822_;
 wire _01823_;
 wire _01824_;
 wire _01825_;
 wire _01826_;
 wire _01827_;
 wire _01828_;
 wire _01829_;
 wire _01830_;
 wire _01831_;
 wire _01832_;
 wire _01833_;
 wire _01834_;
 wire _01835_;
 wire _01836_;
 wire _01837_;
 wire _01838_;
 wire _01839_;
 wire _01840_;
 wire _01841_;
 wire _01842_;
 wire _01843_;
 wire _01844_;
 wire _01845_;
 wire _01846_;
 wire _01847_;
 wire _01848_;
 wire _01849_;
 wire _01850_;
 wire _01851_;
 wire _01852_;
 wire _01853_;
 wire _01854_;
 wire _01855_;
 wire _01856_;
 wire _01857_;
 wire _01858_;
 wire _01859_;
 wire _01860_;
 wire _01861_;
 wire _01862_;
 wire _01863_;
 wire _01864_;
 wire _01865_;
 wire _01866_;
 wire _01867_;
 wire _01868_;
 wire _01869_;
 wire _01870_;
 wire _01871_;
 wire _01872_;
 wire _01873_;
 wire _01874_;
 wire _01875_;
 wire _01876_;
 wire _01877_;
 wire _01878_;
 wire _01879_;
 wire _01880_;
 wire _01881_;
 wire _01882_;
 wire _01883_;
 wire _01884_;
 wire _01885_;
 wire _01886_;
 wire _01887_;
 wire _01888_;
 wire _01889_;
 wire _01890_;
 wire _01891_;
 wire _01892_;
 wire _01893_;
 wire _01894_;
 wire _01895_;
 wire _01896_;
 wire _01897_;
 wire _01898_;
 wire _01899_;
 wire _01900_;
 wire _01901_;
 wire _01902_;
 wire _01903_;
 wire _01904_;
 wire _01905_;
 wire _01906_;
 wire _01907_;
 wire _01908_;
 wire _01909_;
 wire _01910_;
 wire _01911_;
 wire _01912_;
 wire _01913_;
 wire _01914_;
 wire _01915_;
 wire _01916_;
 wire _01917_;
 wire _01918_;
 wire _01919_;
 wire _01920_;
 wire _01921_;
 wire _01922_;
 wire _01923_;
 wire _01924_;
 wire _01925_;
 wire _01926_;
 wire _01927_;
 wire _01928_;
 wire _01929_;
 wire _01930_;
 wire _01931_;
 wire _01932_;
 wire _01933_;
 wire _01934_;
 wire _01935_;
 wire _01936_;
 wire _01937_;
 wire _01938_;
 wire _01939_;
 wire _01940_;
 wire _01941_;
 wire _01942_;
 wire _01943_;
 wire _01944_;
 wire _01945_;
 wire _01946_;
 wire _01947_;
 wire _01948_;
 wire _01949_;
 wire _01950_;
 wire _01951_;
 wire _01952_;
 wire _01953_;
 wire _01954_;
 wire _01955_;
 wire _01956_;
 wire _01957_;
 wire _01958_;
 wire _01959_;
 wire _01960_;
 wire _01961_;
 wire _01962_;
 wire _01963_;
 wire _01964_;
 wire _01965_;
 wire _01966_;
 wire _01967_;
 wire _01968_;
 wire _01969_;
 wire _01970_;
 wire _01971_;
 wire _01972_;
 wire _01973_;
 wire _01974_;
 wire _01975_;
 wire _01976_;
 wire _01977_;
 wire _01978_;
 wire _01979_;
 wire _01980_;
 wire _01981_;
 wire _01982_;
 wire _01983_;
 wire _01984_;
 wire _01985_;
 wire _01986_;
 wire _01987_;
 wire _01988_;
 wire _01989_;
 wire _01990_;
 wire _01991_;
 wire _01992_;
 wire _01993_;
 wire _01994_;
 wire _01995_;
 wire _01996_;
 wire _01997_;
 wire _01998_;
 wire _01999_;
 wire _02000_;
 wire _02001_;
 wire _02002_;
 wire _02003_;
 wire _02004_;
 wire _02005_;
 wire _02006_;
 wire _02007_;
 wire _02008_;
 wire _02009_;
 wire _02010_;
 wire _02011_;
 wire _02012_;
 wire _02013_;
 wire _02014_;
 wire _02015_;
 wire _02016_;
 wire _02017_;
 wire _02018_;
 wire _02019_;
 wire _02020_;
 wire _02021_;
 wire _02022_;
 wire _02023_;
 wire _02024_;
 wire _02025_;
 wire _02026_;
 wire _02027_;
 wire _02028_;
 wire _02029_;
 wire _02030_;
 wire _02031_;
 wire _02032_;
 wire _02033_;
 wire _02034_;
 wire _02035_;
 wire _02036_;
 wire _02037_;
 wire _02038_;
 wire _02039_;
 wire _02040_;
 wire _02041_;
 wire _02042_;
 wire _02043_;
 wire _02044_;
 wire _02045_;
 wire _02046_;
 wire _02047_;
 wire _02048_;
 wire _02049_;
 wire _02050_;
 wire _02051_;
 wire _02052_;
 wire _02053_;
 wire _02054_;
 wire _02055_;
 wire _02056_;
 wire _02057_;
 wire _02058_;
 wire _02059_;
 wire _02060_;
 wire _02061_;
 wire _02062_;
 wire _02063_;
 wire _02064_;
 wire _02065_;
 wire _02066_;
 wire _02067_;
 wire _02068_;
 wire _02069_;
 wire _02070_;
 wire _02071_;
 wire _02072_;
 wire _02073_;
 wire _02074_;
 wire _02075_;
 wire _02076_;
 wire _02077_;
 wire _02078_;
 wire _02079_;
 wire _02080_;
 wire _02081_;
 wire _02082_;
 wire _02083_;
 wire _02084_;
 wire _02085_;
 wire _02086_;
 wire _02087_;
 wire _02088_;
 wire _02089_;
 wire _02090_;
 wire _02091_;
 wire _02092_;
 wire _02093_;
 wire _02094_;
 wire _02095_;
 wire _02096_;
 wire _02097_;
 wire _02098_;
 wire _02099_;
 wire _02100_;
 wire _02101_;
 wire _02102_;
 wire _02103_;
 wire _02104_;
 wire _02105_;
 wire _02106_;
 wire _02107_;
 wire _02108_;
 wire _02109_;
 wire _02110_;
 wire _02111_;
 wire _02112_;
 wire _02113_;
 wire _02114_;
 wire _02115_;
 wire _02116_;
 wire _02117_;
 wire _02118_;
 wire _02119_;
 wire _02120_;
 wire _02121_;
 wire _02122_;
 wire _02123_;
 wire _02124_;
 wire _02125_;
 wire _02126_;
 wire _02127_;
 wire _02128_;
 wire _02129_;
 wire _02130_;
 wire _02131_;
 wire _02132_;
 wire _02133_;
 wire _02134_;
 wire _02135_;
 wire _02136_;
 wire _02137_;
 wire _02138_;
 wire _02139_;
 wire _02140_;
 wire _02141_;
 wire _02142_;
 wire _02143_;
 wire _02144_;
 wire _02145_;
 wire _02146_;
 wire _02147_;
 wire _02148_;
 wire _02149_;
 wire _02150_;
 wire _02151_;
 wire _02152_;
 wire _02153_;
 wire _02154_;
 wire _02155_;
 wire _02156_;
 wire _02157_;
 wire _02158_;
 wire _02159_;
 wire _02160_;
 wire _02161_;
 wire _02162_;
 wire _02163_;
 wire _02164_;
 wire _02165_;
 wire _02166_;
 wire _02167_;
 wire _02168_;
 wire _02169_;
 wire _02170_;
 wire _02171_;
 wire _02172_;
 wire _02173_;
 wire _02174_;
 wire _02175_;
 wire _02176_;
 wire _02177_;
 wire _02178_;
 wire _02179_;
 wire _02180_;
 wire _02181_;
 wire _02182_;
 wire _02183_;
 wire _02184_;
 wire _02185_;
 wire _02186_;
 wire _02187_;
 wire _02188_;
 wire _02189_;
 wire _02190_;
 wire _02191_;
 wire _02192_;
 wire _02193_;
 wire _02194_;
 wire _02195_;
 wire _02196_;
 wire _02197_;
 wire _02198_;
 wire _02199_;
 wire _02200_;
 wire _02201_;
 wire _02202_;
 wire _02203_;
 wire _02204_;
 wire _02205_;
 wire _02206_;
 wire _02207_;
 wire _02208_;
 wire _02209_;
 wire _02210_;
 wire _02211_;
 wire _02212_;
 wire _02213_;
 wire _02214_;
 wire _02215_;
 wire _02216_;
 wire _02217_;
 wire _02218_;
 wire _02219_;
 wire _02220_;
 wire _02221_;
 wire _02222_;
 wire _02223_;
 wire _02224_;
 wire _02225_;
 wire _02226_;
 wire _02227_;
 wire _02228_;
 wire _02229_;
 wire _02230_;
 wire _02231_;
 wire _02232_;
 wire _02233_;
 wire _02234_;
 wire _02235_;
 wire _02236_;
 wire _02237_;
 wire _02238_;
 wire _02239_;
 wire _02240_;
 wire _02241_;
 wire _02242_;
 wire _02243_;
 wire _02244_;
 wire _02245_;
 wire _02246_;
 wire _02247_;
 wire _02248_;
 wire _02249_;
 wire _02250_;
 wire _02251_;
 wire _02252_;
 wire _02253_;
 wire _02254_;
 wire _02255_;
 wire _02256_;
 wire _02257_;
 wire _02258_;
 wire _02259_;
 wire _02260_;
 wire _02261_;
 wire _02262_;
 wire _02263_;
 wire _02264_;
 wire _02265_;
 wire _02266_;
 wire _02267_;
 wire _02268_;
 wire _02269_;
 wire _02270_;
 wire _02271_;
 wire _02272_;
 wire _02273_;
 wire _02274_;
 wire _02275_;
 wire _02276_;
 wire _02277_;
 wire _02278_;
 wire _02279_;
 wire _02280_;
 wire _02281_;
 wire _02282_;
 wire _02283_;
 wire _02284_;
 wire _02285_;
 wire _02286_;
 wire _02287_;
 wire _02288_;
 wire _02289_;
 wire _02290_;
 wire _02291_;
 wire _02292_;
 wire _02293_;
 wire _02294_;
 wire _02295_;
 wire _02296_;
 wire _02297_;
 wire _02298_;
 wire _02299_;
 wire _02300_;
 wire _02301_;
 wire _02302_;
 wire _02303_;
 wire _02304_;
 wire _02305_;
 wire _02306_;
 wire _02307_;
 wire _02308_;
 wire _02309_;
 wire _02310_;
 wire _02311_;
 wire _02312_;
 wire _02313_;
 wire _02314_;
 wire _02315_;
 wire _02316_;
 wire _02317_;
 wire _02318_;
 wire _02319_;
 wire _02320_;
 wire _02321_;
 wire _02322_;
 wire _02323_;
 wire _02324_;
 wire _02325_;
 wire _02326_;
 wire _02327_;
 wire _02328_;
 wire _02329_;
 wire _02330_;
 wire _02331_;
 wire _02332_;
 wire _02333_;
 wire _02334_;
 wire _02335_;
 wire _02336_;
 wire _02337_;
 wire _02338_;
 wire _02339_;
 wire _02340_;
 wire _02341_;
 wire _02342_;
 wire _02343_;
 wire _02344_;
 wire _02345_;
 wire _02346_;
 wire _02347_;
 wire _02348_;
 wire _02349_;
 wire _02350_;
 wire _02351_;
 wire _02352_;
 wire _02353_;
 wire _02354_;
 wire _02355_;
 wire _02356_;
 wire _02357_;
 wire _02358_;
 wire _02359_;
 wire _02360_;
 wire _02361_;
 wire _02362_;
 wire _02363_;
 wire _02364_;
 wire _02365_;
 wire _02366_;
 wire _02367_;
 wire _02368_;
 wire _02369_;
 wire _02370_;
 wire _02371_;
 wire _02372_;
 wire _02373_;
 wire _02374_;
 wire _02375_;
 wire _02376_;
 wire _02377_;
 wire _02378_;
 wire _02379_;
 wire _02380_;
 wire _02381_;
 wire _02382_;
 wire _02383_;
 wire _02384_;
 wire _02385_;
 wire _02386_;
 wire _02387_;
 wire _02388_;
 wire _02389_;
 wire _02390_;
 wire _02391_;
 wire _02392_;
 wire _02393_;
 wire _02394_;
 wire _02395_;
 wire _02396_;
 wire _02397_;
 wire _02398_;
 wire _02399_;
 wire _02400_;
 wire _02401_;
 wire _02402_;
 wire _02403_;
 wire _02404_;
 wire _02405_;
 wire _02406_;
 wire _02407_;
 wire _02408_;
 wire _02409_;
 wire _02410_;
 wire _02411_;
 wire _02412_;
 wire _02413_;
 wire _02414_;
 wire _02415_;
 wire _02416_;
 wire _02417_;
 wire _02418_;
 wire _02419_;
 wire _02420_;
 wire _02421_;
 wire _02422_;
 wire _02423_;
 wire _02424_;
 wire _02425_;
 wire _02426_;
 wire _02427_;
 wire _02428_;
 wire _02429_;
 wire _02430_;
 wire _02431_;
 wire _02432_;
 wire _02433_;
 wire _02434_;
 wire _02435_;
 wire _02436_;
 wire _02437_;
 wire _02438_;
 wire _02439_;
 wire _02440_;
 wire _02441_;
 wire _02442_;
 wire _02443_;
 wire _02444_;
 wire _02445_;
 wire _02446_;
 wire _02447_;
 wire _02448_;
 wire _02449_;
 wire _02450_;
 wire _02451_;
 wire _02452_;
 wire _02453_;
 wire _02454_;
 wire _02455_;
 wire _02456_;
 wire _02457_;
 wire _02458_;
 wire _02459_;
 wire _02460_;
 wire _02461_;
 wire _02462_;
 wire _02463_;
 wire _02464_;
 wire _02465_;
 wire _02466_;
 wire _02467_;
 wire _02468_;
 wire _02469_;
 wire _02470_;
 wire _02471_;
 wire _02472_;
 wire _02473_;
 wire _02474_;
 wire _02475_;
 wire _02476_;
 wire _02477_;
 wire _02478_;
 wire _02479_;
 wire _02480_;
 wire _02481_;
 wire _02482_;
 wire _02483_;
 wire _02484_;
 wire _02485_;
 wire _02486_;
 wire _02487_;
 wire _02488_;
 wire _02489_;
 wire _02490_;
 wire _02491_;
 wire _02492_;
 wire _02493_;
 wire _02494_;
 wire _02495_;
 wire _02496_;
 wire _02497_;
 wire _02498_;
 wire _02499_;
 wire _02500_;
 wire _02501_;
 wire _02502_;
 wire _02503_;
 wire _02504_;
 wire _02505_;
 wire _02506_;
 wire _02507_;
 wire _02508_;
 wire _02509_;
 wire _02510_;
 wire _02511_;
 wire _02512_;
 wire _02513_;
 wire _02514_;
 wire _02515_;
 wire _02516_;
 wire _02517_;
 wire _02518_;
 wire _02519_;
 wire _02520_;
 wire _02521_;
 wire _02522_;
 wire _02523_;
 wire _02524_;
 wire _02525_;
 wire _02526_;
 wire _02527_;
 wire _02528_;
 wire _02529_;
 wire _02530_;
 wire _02531_;
 wire _02532_;
 wire _02533_;
 wire _02534_;
 wire _02535_;
 wire _02536_;
 wire _02537_;
 wire _02538_;
 wire _02539_;
 wire _02540_;
 wire _02541_;
 wire _02542_;
 wire _02543_;
 wire _02544_;
 wire _02545_;
 wire _02546_;
 wire _02547_;
 wire _02548_;
 wire _02549_;
 wire _02550_;
 wire _02551_;
 wire _02552_;
 wire _02553_;
 wire _02554_;
 wire _02555_;
 wire _02556_;
 wire _02557_;
 wire _02558_;
 wire _02559_;
 wire _02560_;
 wire _02561_;
 wire _02562_;
 wire _02563_;
 wire _02564_;
 wire _02565_;
 wire _02566_;
 wire _02567_;
 wire _02568_;
 wire _02569_;
 wire _02570_;
 wire _02571_;
 wire _02572_;
 wire _02573_;
 wire _02574_;
 wire _02575_;
 wire _02576_;
 wire _02577_;
 wire _02578_;
 wire _02579_;
 wire _02580_;
 wire _02581_;
 wire _02582_;
 wire _02583_;
 wire _02584_;
 wire _02585_;
 wire _02586_;
 wire _02587_;
 wire _02588_;
 wire _02589_;
 wire _02590_;
 wire _02591_;
 wire _02592_;
 wire _02593_;
 wire _02594_;
 wire _02595_;
 wire _02596_;
 wire _02597_;
 wire _02598_;
 wire _02599_;
 wire _02600_;
 wire _02601_;
 wire _02602_;
 wire _02603_;
 wire _02604_;
 wire _02605_;
 wire _02606_;
 wire _02607_;
 wire _02608_;
 wire _02609_;
 wire _02610_;
 wire _02611_;
 wire _02612_;
 wire _02613_;
 wire _02614_;
 wire _02615_;
 wire _02616_;
 wire _02617_;
 wire _02618_;
 wire _02619_;
 wire _02620_;
 wire _02621_;
 wire _02622_;
 wire _02623_;
 wire _02624_;
 wire _02625_;
 wire _02626_;
 wire _02627_;
 wire _02628_;
 wire _02629_;
 wire _02630_;
 wire _02631_;
 wire _02632_;
 wire _02633_;
 wire _02634_;
 wire _02635_;
 wire _02636_;
 wire _02637_;
 wire _02638_;
 wire _02639_;
 wire _02640_;
 wire _02641_;
 wire _02642_;
 wire _02643_;
 wire _02644_;
 wire _02645_;
 wire _02646_;
 wire _02647_;
 wire _02648_;
 wire _02649_;
 wire _02650_;
 wire _02651_;
 wire _02652_;
 wire _02653_;
 wire _02654_;
 wire _02655_;
 wire _02656_;
 wire _02657_;
 wire _02658_;
 wire _02659_;
 wire _02660_;
 wire _02661_;
 wire _02662_;
 wire _02663_;
 wire _02664_;
 wire _02665_;
 wire _02666_;
 wire _02667_;
 wire _02668_;
 wire _02669_;
 wire _02670_;
 wire _02671_;
 wire _02672_;
 wire _02673_;
 wire _02674_;
 wire _02675_;
 wire _02676_;
 wire _02677_;
 wire _02678_;
 wire _02679_;
 wire _02680_;
 wire _02681_;
 wire _02682_;
 wire _02683_;
 wire _02684_;
 wire _02685_;
 wire _02686_;
 wire _02687_;
 wire _02688_;
 wire _02689_;
 wire _02690_;
 wire _02691_;
 wire _02692_;
 wire _02693_;
 wire _02694_;
 wire _02695_;
 wire _02696_;
 wire _02697_;
 wire _02698_;
 wire _02699_;
 wire _02700_;
 wire _02701_;
 wire _02702_;
 wire _02703_;
 wire _02704_;
 wire _02705_;
 wire _02706_;
 wire _02707_;
 wire _02708_;
 wire _02709_;
 wire _02710_;
 wire _02711_;
 wire _02712_;
 wire _02713_;
 wire _02714_;
 wire _02715_;
 wire _02716_;
 wire _02717_;
 wire _02718_;
 wire _02719_;
 wire _02720_;
 wire _02721_;
 wire _02722_;
 wire _02723_;
 wire _02724_;
 wire _02725_;
 wire _02726_;
 wire _02727_;
 wire _02728_;
 wire _02729_;
 wire _02730_;
 wire _02731_;
 wire _02732_;
 wire _02733_;
 wire _02734_;
 wire _02735_;
 wire _02736_;
 wire _02737_;
 wire _02738_;
 wire _02739_;
 wire _02740_;
 wire _02741_;
 wire _02742_;
 wire _02743_;
 wire _02744_;
 wire _02745_;
 wire _02746_;
 wire _02747_;
 wire _02748_;
 wire _02749_;
 wire _02750_;
 wire _02751_;
 wire _02752_;
 wire _02753_;
 wire _02754_;
 wire _02755_;
 wire _02756_;
 wire _02757_;
 wire _02758_;
 wire _02759_;
 wire _02760_;
 wire _02761_;
 wire _02762_;
 wire _02763_;
 wire _02764_;
 wire _02765_;
 wire _02766_;
 wire _02767_;
 wire _02768_;
 wire _02769_;
 wire _02770_;
 wire _02771_;
 wire _02772_;
 wire _02773_;
 wire _02774_;
 wire _02775_;
 wire _02776_;
 wire _02777_;
 wire _02778_;
 wire _02779_;
 wire _02780_;
 wire _02781_;
 wire _02782_;
 wire _02783_;
 wire _02784_;
 wire _02785_;
 wire _02786_;
 wire _02787_;
 wire _02788_;
 wire _02789_;
 wire _02790_;
 wire _02791_;
 wire _02792_;
 wire _02793_;
 wire _02794_;
 wire _02795_;
 wire _02796_;
 wire _02797_;
 wire _02798_;
 wire _02799_;
 wire _02800_;
 wire _02801_;
 wire _02802_;
 wire _02803_;
 wire _02804_;
 wire _02805_;
 wire _02806_;
 wire _02807_;
 wire _02808_;
 wire _02809_;
 wire _02810_;
 wire _02811_;
 wire _02812_;
 wire _02813_;
 wire _02814_;
 wire _02815_;
 wire _02816_;
 wire _02817_;
 wire _02818_;
 wire _02819_;
 wire _02820_;
 wire _02821_;
 wire _02822_;
 wire _02823_;
 wire _02824_;
 wire _02825_;
 wire _02826_;
 wire _02827_;
 wire _02828_;
 wire _02829_;
 wire _02830_;
 wire _02831_;
 wire _02832_;
 wire _02833_;
 wire _02834_;
 wire _02835_;
 wire _02836_;
 wire _02837_;
 wire _02838_;
 wire _02839_;
 wire _02840_;
 wire _02841_;
 wire _02842_;
 wire _02843_;
 wire _02844_;
 wire _02845_;
 wire _02846_;
 wire _02847_;
 wire _02848_;
 wire _02849_;
 wire _02850_;
 wire _02851_;
 wire _02852_;
 wire _02853_;
 wire _02854_;
 wire _02855_;
 wire _02856_;
 wire _02857_;
 wire _02858_;
 wire _02859_;
 wire _02860_;
 wire _02861_;
 wire _02862_;
 wire _02863_;
 wire _02864_;
 wire _02865_;
 wire _02866_;
 wire _02867_;
 wire _02868_;
 wire _02869_;
 wire _02870_;
 wire _02871_;
 wire _02872_;
 wire _02873_;
 wire _02874_;
 wire _02875_;
 wire _02876_;
 wire _02877_;
 wire _02878_;
 wire _02879_;
 wire _02880_;
 wire _02881_;
 wire _02882_;
 wire _02883_;
 wire _02884_;
 wire _02885_;
 wire _02886_;
 wire _02887_;
 wire _02888_;
 wire _02889_;
 wire _02890_;
 wire _02891_;
 wire _02892_;
 wire _02893_;
 wire _02894_;
 wire _02895_;
 wire _02896_;
 wire _02897_;
 wire _02898_;
 wire _02899_;
 wire _02900_;
 wire _02901_;
 wire _02902_;
 wire _02903_;
 wire _02904_;
 wire _02905_;
 wire _02906_;
 wire _02907_;
 wire _02908_;
 wire _02909_;
 wire _02910_;
 wire _02911_;
 wire _02912_;
 wire _02913_;
 wire _02914_;
 wire _02915_;
 wire _02916_;
 wire _02917_;
 wire _02918_;
 wire _02919_;
 wire _02920_;
 wire _02921_;
 wire _02922_;
 wire _02923_;
 wire _02924_;
 wire _02925_;
 wire _02926_;
 wire _02927_;
 wire _02928_;
 wire _02929_;
 wire _02930_;
 wire _02931_;
 wire _02932_;
 wire _02933_;
 wire _02934_;
 wire _02935_;
 wire _02936_;
 wire _02937_;
 wire _02938_;
 wire _02939_;
 wire _02940_;
 wire _02941_;
 wire _02942_;
 wire _02943_;
 wire _02944_;
 wire _02945_;
 wire _02946_;
 wire _02947_;
 wire _02948_;
 wire _02949_;
 wire _02950_;
 wire _02951_;
 wire _02952_;
 wire _02953_;
 wire _02954_;
 wire _02955_;
 wire _02956_;
 wire _02957_;
 wire _02958_;
 wire _02959_;
 wire _02960_;
 wire _02961_;
 wire _02962_;
 wire _02963_;
 wire _02964_;
 wire _02965_;
 wire _02966_;
 wire _02967_;
 wire _02968_;
 wire _02969_;
 wire _02970_;
 wire _02971_;
 wire _02972_;
 wire _02973_;
 wire _02974_;
 wire _02975_;
 wire _02976_;
 wire _02977_;
 wire _02978_;
 wire _02979_;
 wire _02980_;
 wire _02981_;
 wire _02982_;
 wire _02983_;
 wire _02984_;
 wire _02985_;
 wire _02986_;
 wire _02987_;
 wire _02988_;
 wire _02989_;
 wire _02990_;
 wire _02991_;
 wire _02992_;
 wire _02993_;
 wire _02994_;
 wire _02995_;
 wire _02996_;
 wire _02997_;
 wire _02998_;
 wire _02999_;
 wire _03000_;
 wire _03001_;
 wire _03002_;
 wire _03003_;
 wire _03004_;
 wire _03005_;
 wire _03006_;
 wire _03007_;
 wire _03008_;
 wire _03009_;
 wire _03010_;
 wire _03011_;
 wire _03012_;
 wire _03013_;
 wire _03014_;
 wire _03015_;
 wire _03016_;
 wire _03017_;
 wire _03018_;
 wire _03019_;
 wire _03020_;
 wire _03021_;
 wire _03022_;
 wire _03023_;
 wire _03024_;
 wire _03025_;
 wire _03026_;
 wire _03027_;
 wire _03028_;
 wire _03029_;
 wire _03030_;
 wire _03031_;
 wire _03032_;
 wire _03033_;
 wire _03034_;
 wire _03035_;
 wire _03036_;
 wire _03037_;
 wire _03038_;
 wire _03039_;
 wire _03040_;
 wire _03041_;
 wire _03042_;
 wire _03043_;
 wire _03044_;
 wire _03045_;
 wire _03046_;
 wire _03047_;
 wire _03048_;
 wire _03049_;
 wire _03050_;
 wire _03051_;
 wire _03052_;
 wire _03053_;
 wire _03054_;
 wire _03055_;
 wire _03056_;
 wire _03057_;
 wire _03058_;
 wire _03059_;
 wire _03060_;
 wire _03061_;
 wire _03062_;
 wire _03063_;
 wire _03064_;
 wire _03065_;
 wire _03066_;
 wire _03067_;
 wire _03068_;
 wire _03069_;
 wire _03070_;
 wire _03071_;
 wire _03072_;
 wire _03073_;
 wire _03074_;
 wire _03075_;
 wire _03076_;
 wire _03077_;
 wire _03078_;
 wire _03079_;
 wire _03080_;
 wire _03081_;
 wire _03082_;
 wire _03083_;
 wire _03084_;
 wire _03085_;
 wire _03086_;
 wire _03087_;
 wire _03088_;
 wire _03089_;
 wire _03090_;
 wire _03091_;
 wire _03092_;
 wire _03093_;
 wire _03094_;
 wire _03095_;
 wire _03096_;
 wire _03097_;
 wire _03098_;
 wire _03099_;
 wire _03100_;
 wire _03101_;
 wire _03102_;
 wire _03103_;
 wire _03104_;
 wire _03105_;
 wire _03106_;
 wire _03107_;
 wire _03108_;
 wire _03109_;
 wire _03110_;
 wire _03111_;
 wire _03112_;
 wire _03113_;
 wire _03114_;
 wire _03115_;
 wire _03116_;
 wire _03117_;
 wire _03118_;
 wire _03119_;
 wire _03120_;
 wire _03121_;
 wire _03122_;
 wire _03123_;
 wire _03124_;
 wire _03125_;
 wire _03126_;
 wire _03127_;
 wire _03128_;
 wire _03129_;
 wire _03130_;
 wire _03131_;
 wire _03132_;
 wire _03133_;
 wire _03134_;
 wire _03135_;
 wire _03136_;
 wire _03137_;
 wire _03138_;
 wire _03139_;
 wire _03140_;
 wire _03141_;
 wire _03142_;
 wire _03143_;
 wire _03144_;
 wire _03145_;
 wire _03146_;
 wire _03147_;
 wire _03148_;
 wire _03149_;
 wire _03150_;
 wire _03151_;
 wire _03152_;
 wire _03153_;
 wire _03154_;
 wire _03155_;
 wire _03156_;
 wire _03157_;
 wire _03158_;
 wire _03159_;
 wire _03160_;
 wire _03161_;
 wire _03162_;
 wire _03163_;
 wire _03164_;
 wire _03165_;
 wire _03166_;
 wire _03167_;
 wire _03168_;
 wire _03169_;
 wire _03170_;
 wire _03171_;
 wire _03172_;
 wire _03173_;
 wire _03174_;
 wire _03175_;
 wire _03176_;
 wire _03177_;
 wire _03178_;
 wire _03179_;
 wire _03180_;
 wire _03181_;
 wire _03182_;
 wire _03183_;
 wire _03184_;
 wire _03185_;
 wire _03186_;
 wire _03187_;
 wire _03188_;
 wire _03189_;
 wire _03190_;
 wire _03191_;
 wire _03192_;
 wire _03193_;
 wire _03194_;
 wire _03195_;
 wire _03196_;
 wire _03197_;
 wire _03198_;
 wire _03199_;
 wire _03200_;
 wire _03201_;
 wire _03202_;
 wire _03203_;
 wire _03204_;
 wire _03205_;
 wire _03206_;
 wire _03207_;
 wire _03208_;
 wire _03209_;
 wire _03210_;
 wire _03211_;
 wire _03212_;
 wire _03213_;
 wire _03214_;
 wire _03215_;
 wire _03216_;
 wire _03217_;
 wire _03218_;
 wire _03219_;
 wire _03220_;
 wire _03221_;
 wire _03222_;
 wire _03223_;
 wire _03224_;
 wire _03225_;
 wire _03226_;
 wire _03227_;
 wire _03228_;
 wire _03229_;
 wire _03230_;
 wire _03231_;
 wire _03232_;
 wire _03233_;
 wire _03234_;
 wire _03235_;
 wire _03236_;
 wire _03237_;
 wire _03238_;
 wire _03239_;
 wire _03240_;
 wire _03241_;
 wire _03242_;
 wire _03243_;
 wire _03244_;
 wire _03245_;
 wire _03246_;
 wire _03247_;
 wire _03248_;
 wire _03249_;
 wire _03250_;
 wire _03251_;
 wire _03252_;
 wire _03253_;
 wire _03254_;
 wire _03255_;
 wire _03256_;
 wire _03257_;
 wire _03258_;
 wire _03259_;
 wire _03260_;
 wire _03261_;
 wire _03262_;
 wire _03263_;
 wire _03264_;
 wire _03265_;
 wire _03266_;
 wire _03267_;
 wire _03268_;
 wire _03269_;
 wire _03270_;
 wire _03271_;
 wire _03272_;
 wire _03273_;
 wire _03274_;
 wire _03275_;
 wire _03276_;
 wire _03277_;
 wire _03278_;
 wire _03279_;
 wire _03280_;
 wire _03281_;
 wire _03282_;
 wire _03283_;
 wire _03284_;
 wire _03285_;
 wire _03286_;
 wire _03287_;
 wire _03288_;
 wire _03289_;
 wire _03290_;
 wire _03291_;
 wire _03292_;
 wire _03293_;
 wire _03294_;
 wire _03295_;
 wire _03296_;
 wire _03297_;
 wire _03298_;
 wire _03299_;
 wire _03300_;
 wire _03301_;
 wire _03302_;
 wire _03303_;
 wire _03304_;
 wire _03305_;
 wire _03306_;
 wire _03307_;
 wire _03308_;
 wire _03309_;
 wire _03310_;
 wire _03311_;
 wire _03312_;
 wire _03313_;
 wire _03314_;
 wire _03315_;
 wire _03316_;
 wire _03317_;
 wire _03318_;
 wire _03319_;
 wire _03320_;
 wire _03321_;
 wire _03322_;
 wire _03323_;
 wire _03324_;
 wire _03325_;
 wire _03326_;
 wire _03327_;
 wire _03328_;
 wire _03329_;
 wire _03330_;
 wire _03331_;
 wire _03332_;
 wire _03333_;
 wire _03334_;
 wire _03335_;
 wire _03336_;
 wire _03337_;
 wire _03338_;
 wire _03339_;
 wire _03340_;
 wire _03341_;
 wire _03342_;
 wire _03343_;
 wire _03344_;
 wire _03345_;
 wire _03346_;
 wire _03347_;
 wire _03348_;
 wire _03349_;
 wire _03350_;
 wire _03351_;
 wire _03352_;
 wire _03353_;
 wire _03354_;
 wire _03355_;
 wire _03356_;
 wire _03357_;
 wire _03358_;
 wire _03359_;
 wire _03360_;
 wire _03361_;
 wire _03362_;
 wire _03363_;
 wire _03364_;
 wire _03365_;
 wire _03366_;
 wire _03367_;
 wire _03368_;
 wire _03369_;
 wire _03370_;
 wire _03371_;
 wire _03372_;
 wire _03373_;
 wire _03374_;
 wire _03375_;
 wire _03376_;
 wire _03377_;
 wire _03378_;
 wire _03379_;
 wire _03380_;
 wire _03381_;
 wire _03382_;
 wire _03383_;
 wire _03384_;
 wire _03385_;
 wire _03386_;
 wire _03387_;
 wire _03388_;
 wire _03389_;
 wire _03390_;
 wire _03391_;
 wire _03392_;
 wire _03393_;
 wire _03394_;
 wire _03395_;
 wire _03396_;
 wire _03397_;
 wire _03398_;
 wire _03399_;
 wire _03400_;
 wire _03401_;
 wire _03402_;
 wire _03403_;
 wire _03404_;
 wire _03405_;
 wire _03406_;
 wire _03407_;
 wire _03408_;
 wire _03409_;
 wire _03410_;
 wire _03411_;
 wire _03412_;
 wire _03413_;
 wire _03414_;
 wire _03415_;
 wire _03416_;
 wire _03417_;
 wire _03418_;
 wire _03419_;
 wire _03420_;
 wire _03421_;
 wire _03422_;
 wire _03423_;
 wire _03424_;
 wire _03425_;
 wire _03426_;
 wire _03427_;
 wire _03428_;
 wire _03429_;
 wire _03430_;
 wire _03431_;
 wire _03432_;
 wire _03433_;
 wire _03434_;
 wire _03435_;
 wire _03436_;
 wire _03437_;
 wire _03438_;
 wire _03439_;
 wire _03440_;
 wire _03441_;
 wire _03442_;
 wire _03443_;
 wire _03444_;
 wire _03445_;
 wire _03446_;
 wire _03447_;
 wire _03448_;
 wire _03449_;
 wire _03450_;
 wire _03451_;
 wire _03452_;
 wire _03453_;
 wire _03454_;
 wire _03455_;
 wire _03456_;
 wire _03457_;
 wire _03458_;
 wire _03459_;
 wire _03460_;
 wire _03461_;
 wire _03462_;
 wire _03463_;
 wire _03464_;
 wire _03465_;
 wire _03466_;
 wire _03467_;
 wire _03468_;
 wire _03469_;
 wire _03470_;
 wire _03471_;
 wire _03472_;
 wire _03473_;
 wire _03474_;
 wire _03475_;
 wire _03476_;
 wire _03477_;
 wire _03478_;
 wire _03479_;
 wire _03480_;
 wire _03481_;
 wire _03482_;
 wire _03483_;
 wire _03484_;
 wire _03485_;
 wire _03486_;
 wire _03487_;
 wire _03488_;
 wire _03489_;
 wire _03490_;
 wire _03491_;
 wire _03492_;
 wire _03493_;
 wire _03494_;
 wire _03495_;
 wire _03496_;
 wire _03497_;
 wire _03498_;
 wire _03499_;
 wire _03500_;
 wire _03501_;
 wire _03502_;
 wire _03503_;
 wire _03504_;
 wire _03505_;
 wire _03506_;
 wire _03507_;
 wire _03508_;
 wire _03509_;
 wire _03510_;
 wire _03511_;
 wire _03512_;
 wire _03513_;
 wire _03514_;
 wire _03515_;
 wire _03516_;
 wire _03517_;
 wire _03518_;
 wire _03519_;
 wire _03520_;
 wire _03521_;
 wire _03522_;
 wire _03523_;
 wire _03524_;
 wire _03525_;
 wire _03526_;
 wire _03527_;
 wire _03528_;
 wire _03529_;
 wire _03530_;
 wire _03531_;
 wire _03532_;
 wire _03533_;
 wire _03534_;
 wire _03535_;
 wire _03536_;
 wire _03537_;
 wire _03538_;
 wire _03539_;
 wire _03540_;
 wire _03541_;
 wire _03542_;
 wire _03543_;
 wire _03544_;
 wire _03545_;
 wire _03546_;
 wire _03547_;
 wire _03548_;
 wire _03549_;
 wire _03550_;
 wire _03551_;
 wire _03552_;
 wire _03553_;
 wire _03554_;
 wire _03555_;
 wire _03556_;
 wire _03557_;
 wire _03558_;
 wire _03559_;
 wire _03560_;
 wire _03561_;
 wire _03562_;
 wire _03563_;
 wire _03564_;
 wire _03565_;
 wire _03566_;
 wire _03567_;
 wire _03568_;
 wire _03569_;
 wire _03570_;
 wire _03571_;
 wire _03572_;
 wire _03573_;
 wire _03574_;
 wire _03575_;
 wire _03576_;
 wire _03577_;
 wire _03578_;
 wire _03579_;
 wire _03580_;
 wire _03581_;
 wire _03582_;
 wire _03583_;
 wire _03584_;
 wire _03585_;
 wire _03586_;
 wire _03587_;
 wire _03588_;
 wire _03589_;
 wire _03590_;
 wire _03591_;
 wire _03592_;
 wire _03593_;
 wire _03594_;
 wire _03595_;
 wire _03596_;
 wire _03597_;
 wire _03598_;
 wire _03599_;
 wire _03600_;
 wire _03601_;
 wire _03602_;
 wire _03603_;
 wire _03604_;
 wire _03605_;
 wire _03606_;
 wire _03607_;
 wire _03608_;
 wire _03609_;
 wire _03610_;
 wire _03611_;
 wire _03612_;
 wire _03613_;
 wire _03614_;
 wire _03615_;
 wire _03616_;
 wire _03617_;
 wire _03618_;
 wire _03619_;
 wire _03620_;
 wire _03621_;
 wire _03622_;
 wire _03623_;
 wire _03624_;
 wire _03625_;
 wire _03626_;
 wire _03627_;
 wire _03628_;
 wire _03629_;
 wire _03630_;
 wire _03631_;
 wire _03632_;
 wire _03633_;
 wire _03634_;
 wire _03635_;
 wire _03636_;
 wire _03637_;
 wire _03638_;
 wire _03639_;
 wire _03640_;
 wire _03641_;
 wire _03642_;
 wire _03643_;
 wire _03644_;
 wire _03645_;
 wire _03646_;
 wire _03647_;
 wire _03648_;
 wire _03649_;
 wire _03650_;
 wire _03651_;
 wire _03652_;
 wire _03653_;
 wire _03654_;
 wire _03655_;
 wire _03656_;
 wire _03657_;
 wire _03658_;
 wire _03659_;
 wire _03660_;
 wire _03661_;
 wire _03662_;
 wire _03663_;
 wire _03664_;
 wire _03665_;
 wire _03666_;
 wire _03667_;
 wire _03668_;
 wire _03669_;
 wire _03670_;
 wire _03671_;
 wire _03672_;
 wire _03673_;
 wire _03674_;
 wire _03675_;
 wire _03676_;
 wire _03677_;
 wire _03678_;
 wire _03679_;
 wire _03680_;
 wire _03681_;
 wire _03682_;
 wire _03683_;
 wire _03684_;
 wire _03685_;
 wire _03686_;
 wire _03687_;
 wire _03688_;
 wire _03689_;
 wire _03690_;
 wire _03691_;
 wire _03692_;
 wire _03693_;
 wire _03694_;
 wire _03695_;
 wire _03696_;
 wire _03697_;
 wire _03698_;
 wire _03699_;
 wire _03700_;
 wire _03701_;
 wire _03702_;
 wire _03703_;
 wire _03704_;
 wire _03705_;
 wire _03706_;
 wire _03707_;
 wire _03708_;
 wire _03709_;
 wire _03710_;
 wire _03711_;
 wire _03712_;
 wire _03713_;
 wire _03714_;
 wire _03715_;
 wire _03716_;
 wire _03717_;
 wire _03718_;
 wire _03719_;
 wire _03720_;
 wire _03721_;
 wire _03722_;
 wire _03723_;
 wire _03724_;
 wire _03725_;
 wire _03726_;
 wire _03727_;
 wire _03728_;
 wire _03729_;
 wire _03730_;
 wire _03731_;
 wire _03732_;
 wire _03733_;
 wire _03734_;
 wire _03735_;
 wire _03736_;
 wire _03737_;
 wire _03738_;
 wire _03739_;
 wire _03740_;
 wire _03741_;
 wire _03742_;
 wire _03743_;
 wire _03744_;
 wire _03745_;
 wire _03746_;
 wire _03747_;
 wire _03748_;
 wire _03749_;
 wire _03750_;
 wire _03751_;
 wire _03752_;
 wire _03753_;
 wire _03754_;
 wire _03755_;
 wire _03756_;
 wire _03757_;
 wire _03758_;
 wire _03759_;
 wire _03760_;
 wire _03761_;
 wire _03762_;
 wire _03763_;
 wire _03764_;
 wire _03765_;
 wire _03766_;
 wire _03767_;
 wire _03768_;
 wire _03769_;
 wire _03770_;
 wire _03771_;
 wire _03772_;
 wire _03773_;
 wire _03774_;
 wire _03775_;
 wire _03776_;
 wire _03777_;
 wire _03778_;
 wire _03779_;
 wire _03780_;
 wire _03781_;
 wire _03782_;
 wire _03783_;
 wire _03784_;
 wire _03785_;
 wire _03786_;
 wire _03787_;
 wire _03788_;
 wire _03789_;
 wire _03790_;
 wire _03791_;
 wire _03792_;
 wire _03793_;
 wire _03794_;
 wire _03795_;
 wire _03796_;
 wire _03797_;
 wire _03798_;
 wire _03799_;
 wire _03800_;
 wire _03801_;
 wire _03802_;
 wire _03803_;
 wire _03804_;
 wire _03805_;
 wire _03806_;
 wire _03807_;
 wire _03808_;
 wire _03809_;
 wire _03810_;
 wire _03811_;
 wire _03812_;
 wire _03813_;
 wire _03814_;
 wire _03815_;
 wire _03816_;
 wire _03817_;
 wire _03818_;
 wire _03819_;
 wire _03820_;
 wire _03821_;
 wire _03822_;
 wire _03823_;
 wire _03824_;
 wire _03825_;
 wire _03826_;
 wire _03827_;
 wire _03828_;
 wire _03829_;
 wire _03830_;
 wire _03831_;
 wire _03832_;
 wire _03833_;
 wire _03834_;
 wire _03835_;
 wire _03836_;
 wire _03837_;
 wire _03838_;
 wire _03839_;
 wire _03840_;
 wire _03841_;
 wire _03842_;
 wire _03843_;
 wire _03844_;
 wire _03845_;
 wire _03846_;
 wire _03847_;
 wire _03848_;
 wire _03849_;
 wire _03850_;
 wire _03851_;
 wire _03852_;
 wire _03853_;
 wire _03854_;
 wire _03855_;
 wire _03856_;
 wire _03857_;
 wire _03858_;
 wire _03859_;
 wire _03860_;
 wire _03861_;
 wire _03862_;
 wire _03863_;
 wire _03864_;
 wire _03865_;
 wire _03866_;
 wire _03867_;
 wire _03868_;
 wire _03869_;
 wire _03870_;
 wire _03871_;
 wire _03872_;
 wire _03873_;
 wire _03874_;
 wire _03875_;
 wire _03876_;
 wire _03877_;
 wire _03878_;
 wire _03879_;
 wire _03880_;
 wire _03881_;
 wire _03882_;
 wire _03883_;
 wire _03884_;
 wire _03885_;
 wire _03886_;
 wire _03887_;
 wire _03888_;
 wire _03889_;
 wire _03890_;
 wire _03891_;
 wire _03892_;
 wire _03893_;
 wire _03894_;
 wire _03895_;
 wire _03896_;
 wire _03897_;
 wire _03898_;
 wire _03899_;
 wire _03900_;
 wire _03901_;
 wire _03902_;
 wire _03903_;
 wire _03904_;
 wire _03905_;
 wire _03906_;
 wire _03907_;
 wire _03908_;
 wire _03909_;
 wire _03910_;
 wire _03911_;
 wire _03912_;
 wire _03913_;
 wire _03914_;
 wire _03915_;
 wire _03916_;
 wire _03917_;
 wire _03918_;
 wire _03919_;
 wire _03920_;
 wire _03921_;
 wire _03922_;
 wire _03923_;
 wire _03924_;
 wire _03925_;
 wire _03926_;
 wire _03927_;
 wire _03928_;
 wire _03929_;
 wire _03930_;
 wire _03931_;
 wire _03932_;
 wire _03933_;
 wire _03934_;
 wire _03935_;
 wire _03936_;
 wire _03937_;
 wire _03938_;
 wire _03939_;
 wire _03940_;
 wire _03941_;
 wire _03942_;
 wire _03943_;
 wire _03944_;
 wire _03945_;
 wire _03946_;
 wire _03947_;
 wire _03948_;
 wire _03949_;
 wire _03950_;
 wire _03951_;
 wire _03952_;
 wire _03953_;
 wire _03954_;
 wire _03955_;
 wire _03956_;
 wire _03957_;
 wire _03958_;
 wire _03959_;
 wire _03960_;
 wire _03961_;
 wire _03962_;
 wire _03963_;
 wire _03964_;
 wire _03965_;
 wire _03966_;
 wire _03967_;
 wire _03968_;
 wire _03969_;
 wire _03970_;
 wire _03971_;
 wire _03972_;
 wire _03973_;
 wire _03974_;
 wire _03975_;
 wire _03976_;
 wire _03977_;
 wire _03978_;
 wire _03979_;
 wire _03980_;
 wire _03981_;
 wire _03982_;
 wire _03983_;
 wire _03984_;
 wire _03985_;
 wire _03986_;
 wire _03987_;
 wire _03988_;
 wire _03989_;
 wire _03990_;
 wire _03991_;
 wire _03992_;
 wire _03993_;
 wire _03994_;
 wire _03995_;
 wire _03996_;
 wire _03997_;
 wire _03998_;
 wire _03999_;
 wire _04000_;
 wire _04001_;
 wire _04002_;
 wire _04003_;
 wire _04004_;
 wire _04005_;
 wire _04006_;
 wire _04007_;
 wire _04008_;
 wire _04009_;
 wire _04010_;
 wire _04011_;
 wire _04012_;
 wire _04013_;
 wire _04014_;
 wire _04015_;
 wire _04016_;
 wire _04017_;
 wire _04018_;
 wire _04019_;
 wire _04020_;
 wire _04021_;
 wire _04022_;
 wire _04023_;
 wire _04024_;
 wire _04025_;
 wire _04026_;
 wire _04027_;
 wire _04028_;
 wire _04029_;
 wire _04030_;
 wire _04031_;
 wire _04032_;
 wire _04033_;
 wire _04034_;
 wire _04035_;
 wire _04036_;
 wire _04037_;
 wire _04038_;
 wire _04039_;
 wire _04040_;
 wire _04041_;
 wire _04042_;
 wire _04043_;
 wire _04044_;
 wire _04045_;
 wire _04046_;
 wire _04047_;
 wire _04048_;
 wire _04049_;
 wire _04050_;
 wire _04051_;
 wire _04052_;
 wire _04053_;
 wire _04054_;
 wire _04055_;
 wire _04056_;
 wire _04057_;
 wire _04058_;
 wire _04059_;
 wire _04060_;
 wire _04061_;
 wire _04062_;
 wire _04063_;
 wire _04064_;
 wire _04065_;
 wire _04066_;
 wire _04067_;
 wire _04068_;
 wire _04069_;
 wire _04070_;
 wire _04071_;
 wire _04072_;
 wire _04073_;
 wire _04074_;
 wire _04075_;
 wire _04076_;
 wire _04077_;
 wire _04078_;
 wire _04079_;
 wire _04080_;
 wire _04081_;
 wire _04082_;
 wire _04083_;
 wire _04084_;
 wire _04085_;
 wire _04086_;
 wire _04087_;
 wire _04088_;
 wire _04089_;
 wire _04090_;
 wire _04091_;
 wire _04092_;
 wire _04093_;
 wire _04094_;
 wire _04095_;
 wire _04096_;
 wire _04097_;
 wire _04098_;
 wire _04099_;
 wire _04100_;
 wire _04101_;
 wire _04102_;
 wire _04103_;
 wire _04104_;
 wire _04105_;
 wire _04106_;
 wire _04107_;
 wire _04108_;
 wire _04109_;
 wire _04110_;
 wire _04111_;
 wire _04112_;
 wire _04113_;
 wire _04114_;
 wire _04115_;
 wire _04116_;
 wire _04117_;
 wire _04118_;
 wire _04119_;
 wire _04120_;
 wire _04121_;
 wire _04122_;
 wire _04123_;
 wire _04124_;
 wire _04125_;
 wire _04126_;
 wire _04127_;
 wire _04128_;
 wire _04129_;
 wire _04130_;
 wire _04131_;
 wire _04132_;
 wire _04133_;
 wire _04134_;
 wire _04135_;
 wire _04136_;
 wire _04137_;
 wire _04138_;
 wire _04139_;
 wire _04140_;
 wire _04141_;
 wire _04142_;
 wire _04143_;
 wire _04144_;
 wire _04145_;
 wire _04146_;
 wire _04147_;
 wire _04148_;
 wire _04149_;
 wire _04150_;
 wire _04151_;
 wire _04152_;
 wire _04153_;
 wire _04154_;
 wire _04155_;
 wire _04156_;
 wire _04157_;
 wire _04158_;
 wire _04159_;
 wire _04160_;
 wire _04161_;
 wire _04162_;
 wire _04163_;
 wire _04164_;
 wire _04165_;
 wire _04166_;
 wire _04167_;
 wire _04168_;
 wire _04169_;
 wire _04170_;
 wire _04171_;
 wire _04172_;
 wire _04173_;
 wire _04174_;
 wire _04175_;
 wire _04176_;
 wire _04177_;
 wire _04178_;
 wire _04179_;
 wire _04180_;
 wire _04181_;
 wire _04182_;
 wire _04183_;
 wire _04184_;
 wire _04185_;
 wire _04186_;
 wire _04187_;
 wire _04188_;
 wire _04189_;
 wire _04190_;
 wire _04191_;
 wire _04192_;
 wire _04193_;
 wire _04194_;
 wire _04195_;
 wire _04196_;
 wire _04197_;
 wire _04198_;
 wire _04199_;
 wire _04200_;
 wire _04201_;
 wire _04202_;
 wire _04203_;
 wire _04204_;
 wire _04205_;
 wire _04206_;
 wire _04207_;
 wire _04208_;
 wire _04209_;
 wire _04210_;
 wire _04211_;
 wire _04212_;
 wire _04213_;
 wire _04214_;
 wire _04215_;
 wire _04216_;
 wire _04217_;
 wire _04218_;
 wire _04219_;
 wire _04220_;
 wire _04221_;
 wire _04222_;
 wire _04223_;
 wire _04224_;
 wire _04225_;
 wire _04226_;
 wire _04227_;
 wire _04228_;
 wire _04229_;
 wire _04230_;
 wire _04231_;
 wire _04232_;
 wire _04233_;
 wire _04234_;
 wire _04235_;
 wire _04236_;
 wire _04237_;
 wire _04238_;
 wire _04239_;
 wire _04240_;
 wire _04241_;
 wire _04242_;
 wire _04243_;
 wire _04244_;
 wire _04245_;
 wire _04246_;
 wire _04247_;
 wire _04248_;
 wire _04249_;
 wire _04250_;
 wire _04251_;
 wire _04252_;
 wire _04253_;
 wire _04254_;
 wire _04255_;
 wire _04256_;
 wire _04257_;
 wire _04258_;
 wire _04259_;
 wire _04260_;
 wire _04261_;
 wire _04262_;
 wire _04263_;
 wire _04264_;
 wire _04265_;
 wire _04266_;
 wire _04267_;
 wire _04268_;
 wire _04269_;
 wire _04270_;
 wire _04271_;
 wire _04272_;
 wire _04273_;
 wire _04274_;
 wire _04275_;
 wire _04276_;
 wire _04277_;
 wire _04278_;
 wire _04279_;
 wire _04280_;
 wire _04281_;
 wire _04282_;
 wire _04283_;
 wire _04284_;
 wire _04285_;
 wire _04286_;
 wire _04287_;
 wire _04288_;
 wire _04289_;
 wire _04290_;
 wire _04291_;
 wire _04292_;
 wire _04293_;
 wire _04294_;
 wire _04295_;
 wire _04296_;
 wire _04297_;
 wire _04298_;
 wire _04299_;
 wire _04300_;
 wire _04301_;
 wire _04302_;
 wire _04303_;
 wire _04304_;
 wire _04305_;
 wire _04306_;
 wire _04307_;
 wire _04308_;
 wire _04309_;
 wire _04310_;
 wire _04311_;
 wire _04312_;
 wire _04313_;
 wire _04314_;
 wire _04315_;
 wire _04316_;
 wire _04317_;
 wire _04318_;
 wire _04319_;
 wire _04320_;
 wire _04321_;
 wire _04322_;
 wire _04323_;
 wire _04324_;
 wire _04325_;
 wire _04326_;
 wire _04327_;
 wire _04328_;
 wire _04329_;
 wire _04330_;
 wire _04331_;
 wire _04332_;
 wire _04333_;
 wire _04334_;
 wire _04335_;
 wire _04336_;
 wire _04337_;
 wire _04338_;
 wire _04339_;
 wire _04340_;
 wire _04341_;
 wire _04342_;
 wire _04343_;
 wire _04344_;
 wire _04345_;
 wire _04346_;
 wire _04347_;
 wire _04353_;
 wire _04354_;
 wire _04355_;
 wire _04356_;
 wire _04357_;
 wire _04358_;
 wire _04359_;
 wire _04360_;
 wire _04361_;
 wire _04362_;
 wire _04363_;
 wire _04364_;
 wire _04365_;
 wire _04366_;
 wire _04367_;
 wire _04368_;
 wire _04369_;
 wire _04370_;
 wire _04371_;
 wire _04372_;
 wire _04373_;
 wire _04374_;
 wire _04375_;
 wire _04376_;
 wire _04377_;
 wire _04378_;
 wire _04379_;
 wire _04380_;
 wire _04381_;
 wire _04382_;
 wire _04383_;
 wire _04384_;
 wire _04385_;
 wire _04386_;
 wire _04387_;
 wire _04388_;
 wire _04389_;
 wire _04390_;
 wire _04391_;
 wire _04392_;
 wire _04393_;
 wire _04394_;
 wire _04395_;
 wire _04396_;
 wire _04397_;
 wire _04398_;
 wire _04399_;
 wire _04400_;
 wire _04401_;
 wire _04402_;
 wire _04403_;
 wire _04404_;
 wire _04405_;
 wire _04406_;
 wire _04407_;
 wire _04408_;
 wire _04409_;
 wire _04410_;
 wire _04411_;
 wire _04412_;
 wire _04413_;
 wire _04414_;
 wire _04415_;
 wire _04416_;
 wire _04417_;
 wire _04418_;
 wire _04419_;
 wire _04420_;
 wire _04421_;
 wire _04422_;
 wire _04423_;
 wire _04424_;
 wire _04425_;
 wire _04426_;
 wire _04427_;
 wire _04428_;
 wire _04429_;
 wire _04430_;
 wire _04431_;
 wire _04432_;
 wire _04433_;
 wire _04434_;
 wire _04435_;
 wire _04436_;
 wire _04437_;
 wire _04438_;
 wire _04439_;
 wire _04440_;
 wire _04441_;
 wire _04442_;
 wire _04443_;
 wire _04444_;
 wire _04445_;
 wire _04446_;
 wire _04447_;
 wire _04448_;
 wire _04449_;
 wire _04450_;
 wire _04451_;
 wire _04452_;
 wire _04453_;
 wire _04454_;
 wire _04455_;
 wire _04456_;
 wire _04457_;
 wire _04458_;
 wire _04459_;
 wire _04460_;
 wire _04461_;
 wire _04462_;
 wire _04463_;
 wire _04464_;
 wire _04465_;
 wire _04466_;
 wire _04467_;
 wire _04468_;
 wire _04469_;
 wire _04470_;
 wire _04471_;
 wire _04472_;
 wire _04473_;
 wire _04474_;
 wire _04475_;
 wire _04476_;
 wire _04477_;
 wire _04478_;
 wire _04479_;
 wire _04480_;
 wire _04481_;
 wire _04482_;
 wire _04483_;
 wire _04484_;
 wire _04485_;
 wire _04486_;
 wire _04487_;
 wire _04488_;
 wire _04489_;
 wire _04490_;
 wire _04491_;
 wire _04492_;
 wire _04493_;
 wire _04494_;
 wire _04495_;
 wire _04496_;
 wire _04497_;
 wire _04498_;
 wire _04499_;
 wire _04500_;
 wire _04501_;
 wire _04502_;
 wire _04503_;
 wire _04504_;
 wire _04505_;
 wire _04506_;
 wire _04507_;
 wire _04508_;
 wire _04509_;
 wire _04510_;
 wire _04511_;
 wire _04512_;
 wire _04513_;
 wire _04514_;
 wire _04515_;
 wire _04516_;
 wire _04517_;
 wire _04518_;
 wire _04519_;
 wire _04520_;
 wire _04521_;
 wire _04522_;
 wire _04523_;
 wire _04524_;
 wire _04525_;
 wire _04526_;
 wire _04527_;
 wire _04528_;
 wire _04529_;
 wire _04530_;
 wire _04531_;
 wire _04532_;
 wire _04533_;
 wire _04534_;
 wire _04535_;
 wire _04536_;
 wire _04537_;
 wire _04538_;
 wire _04539_;
 wire _04540_;
 wire _04541_;
 wire _04542_;
 wire _04543_;
 wire _04544_;
 wire _04545_;
 wire _04546_;
 wire _04547_;
 wire _04548_;
 wire _04549_;
 wire _04550_;
 wire _04551_;
 wire _04552_;
 wire _04553_;
 wire _04554_;
 wire _04555_;
 wire _04556_;
 wire _04557_;
 wire _04558_;
 wire _04559_;
 wire _04560_;
 wire _04561_;
 wire _04562_;
 wire _04563_;
 wire _04564_;
 wire _04565_;
 wire _04566_;
 wire _04567_;
 wire _04568_;
 wire _04569_;
 wire _04570_;
 wire _04571_;
 wire _04572_;
 wire _04573_;
 wire _04574_;
 wire _04575_;
 wire _04576_;
 wire _04577_;
 wire _04578_;
 wire _04579_;
 wire _04580_;
 wire _04581_;
 wire _04582_;
 wire _04583_;
 wire _04584_;
 wire _04585_;
 wire _04586_;
 wire _04587_;
 wire _04588_;
 wire _04589_;
 wire _04590_;
 wire _04591_;
 wire _04592_;
 wire _04593_;
 wire _04594_;
 wire _04595_;
 wire _04596_;
 wire _04597_;
 wire _04598_;
 wire _04599_;
 wire _04600_;
 wire _04601_;
 wire _04602_;
 wire _04603_;
 wire _04604_;
 wire _04605_;
 wire _04606_;
 wire _04607_;
 wire _04608_;
 wire _04609_;
 wire _04610_;
 wire _04611_;
 wire _04612_;
 wire _04613_;
 wire _04614_;
 wire _04615_;
 wire _04616_;
 wire _04617_;
 wire _04618_;
 wire _04619_;
 wire _04620_;
 wire _04621_;
 wire _04622_;
 wire _04623_;
 wire _04624_;
 wire _04625_;
 wire _04626_;
 wire _04627_;
 wire _04628_;
 wire _04629_;
 wire _04630_;
 wire _04631_;
 wire _04632_;
 wire _04633_;
 wire _04634_;
 wire _04635_;
 wire _04636_;
 wire _04637_;
 wire _04638_;
 wire _04639_;
 wire _04640_;
 wire _04641_;
 wire _04642_;
 wire _04643_;
 wire _04644_;
 wire _04645_;
 wire _04646_;
 wire _04647_;
 wire _04648_;
 wire _04649_;
 wire _04650_;
 wire _04651_;
 wire _04652_;
 wire _04653_;
 wire _04654_;
 wire _04655_;
 wire _04656_;
 wire _04657_;
 wire _04658_;
 wire _04659_;
 wire _04660_;
 wire _04661_;
 wire _04662_;
 wire _04663_;
 wire _04664_;
 wire _04665_;
 wire _04666_;
 wire _04667_;
 wire _04668_;
 wire _04669_;
 wire _04670_;
 wire _04671_;
 wire _04672_;
 wire _04673_;
 wire _04674_;
 wire _04675_;
 wire _04676_;
 wire _04677_;
 wire _04678_;
 wire _04679_;
 wire _04680_;
 wire _04681_;
 wire _04682_;
 wire _04683_;
 wire _04684_;
 wire _04685_;
 wire _04686_;
 wire _04687_;
 wire clknet_0__04347_;
 wire clknet_0__04353_;
 wire clknet_0__04354_;
 wire clknet_0__04355_;
 wire clknet_0__04356_;
 wire clknet_0__04357_;
 wire clknet_0__04358_;
 wire clknet_0__04359_;
 wire clknet_0__04392_;
 wire clknet_0__04393_;
 wire clknet_0__04394_;
 wire clknet_0__04395_;
 wire clknet_0__04396_;
 wire clknet_0__04397_;
 wire clknet_0__04398_;
 wire clknet_0__04399_;
 wire clknet_0__04400_;
 wire clknet_0__04401_;
 wire clknet_0__04402_;
 wire clknet_0__04403_;
 wire clknet_0__04404_;
 wire clknet_0__04405_;
 wire clknet_0__04406_;
 wire clknet_0__04407_;
 wire clknet_0__04408_;
 wire clknet_0__04409_;
 wire clknet_0__04410_;
 wire clknet_0__04411_;
 wire clknet_0__04412_;
 wire clknet_0__04413_;
 wire clknet_0__04414_;
 wire clknet_0__04415_;
 wire clknet_0__04416_;
 wire clknet_0__04417_;
 wire clknet_0__04418_;
 wire clknet_0__04419_;
 wire clknet_0__04420_;
 wire clknet_0__04421_;
 wire clknet_0__04422_;
 wire clknet_0__04423_;
 wire clknet_0__04424_;
 wire clknet_0__04425_;
 wire clknet_0__04426_;
 wire clknet_0__04427_;
 wire clknet_0__04428_;
 wire clknet_0__04429_;
 wire clknet_0__04430_;
 wire clknet_0__04431_;
 wire clknet_0__04432_;
 wire clknet_0__04433_;
 wire clknet_0__04434_;
 wire clknet_0__04435_;
 wire clknet_0__04436_;
 wire clknet_0__04437_;
 wire clknet_0__04438_;
 wire clknet_0__04439_;
 wire clknet_0__04440_;
 wire clknet_0__04441_;
 wire clknet_0__04442_;
 wire clknet_0__04443_;
 wire clknet_0__04444_;
 wire clknet_0__04445_;
 wire clknet_0__04446_;
 wire clknet_0__04447_;
 wire clknet_0__04448_;
 wire clknet_0__04449_;
 wire clknet_0__04450_;
 wire clknet_0__04451_;
 wire clknet_0__04452_;
 wire clknet_0__04453_;
 wire clknet_0__04454_;
 wire clknet_0__04455_;
 wire clknet_0__04456_;
 wire clknet_0__04457_;
 wire clknet_0__04458_;
 wire clknet_0__04459_;
 wire clknet_0__04460_;
 wire clknet_0__04461_;
 wire clknet_0__04463_;
 wire clknet_0__04464_;
 wire clknet_0__04465_;
 wire clknet_0__04466_;
 wire clknet_0__04467_;
 wire clknet_0__04468_;
 wire clknet_0__04469_;
 wire clknet_0__04470_;
 wire clknet_0__04471_;
 wire clknet_0__04472_;
 wire clknet_0__04473_;
 wire clknet_0__04474_;
 wire clknet_0__04475_;
 wire clknet_0__04476_;
 wire clknet_0__04477_;
 wire clknet_0__04478_;
 wire clknet_0__04479_;
 wire clknet_0__04480_;
 wire clknet_0__04481_;
 wire clknet_0__04482_;
 wire clknet_0__04483_;
 wire clknet_0__04484_;
 wire clknet_0__04485_;
 wire clknet_0__04486_;
 wire clknet_0__04487_;
 wire clknet_0__04488_;
 wire clknet_0__04489_;
 wire clknet_0__04490_;
 wire clknet_0__04491_;
 wire clknet_0__04492_;
 wire clknet_0__04493_;
 wire clknet_0__04494_;
 wire clknet_0__04495_;
 wire clknet_0__04496_;
 wire clknet_0__04497_;
 wire clknet_0__04498_;
 wire clknet_0__04499_;
 wire clknet_0__04500_;
 wire clknet_0__04501_;
 wire clknet_0__04502_;
 wire clknet_0__04503_;
 wire clknet_0__04504_;
 wire clknet_0__04505_;
 wire clknet_0__04538_;
 wire clknet_0__04539_;
 wire clknet_0__04540_;
 wire clknet_0__04541_;
 wire clknet_0__04542_;
 wire clknet_0__04543_;
 wire clknet_0__04544_;
 wire clknet_0__04545_;
 wire clknet_0__04546_;
 wire clknet_0__04547_;
 wire clknet_0__04548_;
 wire clknet_0__04549_;
 wire clknet_0__04550_;
 wire clknet_0__04551_;
 wire clknet_0__04552_;
 wire clknet_0__04562_;
 wire clknet_0__04564_;
 wire clknet_0__04565_;
 wire clknet_0__04566_;
 wire clknet_0__04567_;
 wire clknet_0__04568_;
 wire clknet_0__04569_;
 wire clknet_0__04570_;
 wire clknet_0__04571_;
 wire clknet_0__04572_;
 wire clknet_0__04573_;
 wire clknet_0__04574_;
 wire clknet_0__04575_;
 wire clknet_0__04576_;
 wire clknet_0__04577_;
 wire clknet_0__04578_;
 wire clknet_0__04579_;
 wire clknet_0__04580_;
 wire clknet_0__04581_;
 wire clknet_0__04582_;
 wire clknet_0__04583_;
 wire clknet_0__04584_;
 wire clknet_0__04586_;
 wire clknet_0__04587_;
 wire clknet_0__04588_;
 wire clknet_0__04589_;
 wire clknet_0__04590_;
 wire clknet_0__04591_;
 wire clknet_0__04592_;
 wire clknet_0__04593_;
 wire clknet_0__04594_;
 wire clknet_0__04595_;
 wire clknet_0__04596_;
 wire clknet_0__04597_;
 wire clknet_0__04598_;
 wire clknet_0__04599_;
 wire clknet_0__04600_;
 wire clknet_0__04601_;
 wire clknet_0__04602_;
 wire clknet_0__04603_;
 wire clknet_0__04604_;
 wire clknet_0__04605_;
 wire clknet_0__04606_;
 wire clknet_0__04608_;
 wire clknet_0__04609_;
 wire clknet_0__04610_;
 wire clknet_0__04611_;
 wire clknet_0__04612_;
 wire clknet_0__04613_;
 wire clknet_0__04614_;
 wire clknet_0__04615_;
 wire clknet_0__04616_;
 wire clknet_0__04617_;
 wire clknet_0__04618_;
 wire clknet_0__04619_;
 wire clknet_0__04620_;
 wire clknet_0__04621_;
 wire clknet_0__04622_;
 wire clknet_0__04623_;
 wire clknet_0__04624_;
 wire clknet_0__04625_;
 wire clknet_0__04626_;
 wire clknet_0__04627_;
 wire clknet_0__04628_;
 wire clknet_0__04629_;
 wire clknet_0__04630_;
 wire clknet_0__04631_;
 wire clknet_0__04632_;
 wire clknet_0__04633_;
 wire clknet_0__04634_;
 wire clknet_0__04635_;
 wire clknet_0__04636_;
 wire clknet_0__04637_;
 wire clknet_0__04638_;
 wire clknet_0__04639_;
 wire clknet_0__04640_;
 wire clknet_0__04641_;
 wire clknet_0__04642_;
 wire clknet_0__04643_;
 wire clknet_0__04644_;
 wire clknet_0__04645_;
 wire clknet_0__04646_;
 wire clknet_0__04647_;
 wire clknet_0__04648_;
 wire clknet_0__04649_;
 wire clknet_0__04650_;
 wire clknet_0__04651_;
 wire clknet_0__04652_;
 wire clknet_0__04653_;
 wire clknet_0__04658_;
 wire clknet_0__04659_;
 wire clknet_0__04664_;
 wire clknet_0__04665_;
 wire clknet_0__04670_;
 wire clknet_0__04671_;
 wire clknet_0__04672_;
 wire clknet_0__04673_;
 wire clknet_0__04674_;
 wire clknet_0__04675_;
 wire clknet_0__04676_;
 wire clknet_0__04679_;
 wire clknet_0__04680_;
 wire clknet_0__04682_;
 wire clknet_0__04685_;
 wire clknet_0__04686_;
 wire clknet_0_mclk;
 wire clknet_0_user_clock1;
 wire clknet_0_user_clock2;
 wire clknet_1_0__leaf__04347_;
 wire clknet_1_0__leaf__04354_;
 wire clknet_1_0__leaf__04355_;
 wire clknet_1_0__leaf__04356_;
 wire clknet_1_0__leaf__04357_;
 wire clknet_1_0__leaf__04392_;
 wire clknet_1_0__leaf__04393_;
 wire clknet_1_0__leaf__04394_;
 wire clknet_1_0__leaf__04395_;
 wire clknet_1_0__leaf__04396_;
 wire clknet_1_0__leaf__04397_;
 wire clknet_1_0__leaf__04398_;
 wire clknet_1_0__leaf__04399_;
 wire clknet_1_0__leaf__04400_;
 wire clknet_1_0__leaf__04401_;
 wire clknet_1_0__leaf__04402_;
 wire clknet_1_0__leaf__04403_;
 wire clknet_1_0__leaf__04404_;
 wire clknet_1_0__leaf__04405_;
 wire clknet_1_0__leaf__04406_;
 wire clknet_1_0__leaf__04407_;
 wire clknet_1_0__leaf__04408_;
 wire clknet_1_0__leaf__04409_;
 wire clknet_1_0__leaf__04410_;
 wire clknet_1_0__leaf__04411_;
 wire clknet_1_0__leaf__04412_;
 wire clknet_1_0__leaf__04413_;
 wire clknet_1_0__leaf__04414_;
 wire clknet_1_0__leaf__04415_;
 wire clknet_1_0__leaf__04416_;
 wire clknet_1_0__leaf__04417_;
 wire clknet_1_0__leaf__04418_;
 wire clknet_1_0__leaf__04419_;
 wire clknet_1_0__leaf__04420_;
 wire clknet_1_0__leaf__04421_;
 wire clknet_1_0__leaf__04422_;
 wire clknet_1_0__leaf__04423_;
 wire clknet_1_0__leaf__04424_;
 wire clknet_1_0__leaf__04425_;
 wire clknet_1_0__leaf__04426_;
 wire clknet_1_0__leaf__04427_;
 wire clknet_1_0__leaf__04428_;
 wire clknet_1_0__leaf__04429_;
 wire clknet_1_0__leaf__04430_;
 wire clknet_1_0__leaf__04431_;
 wire clknet_1_0__leaf__04432_;
 wire clknet_1_0__leaf__04433_;
 wire clknet_1_0__leaf__04434_;
 wire clknet_1_0__leaf__04435_;
 wire clknet_1_0__leaf__04436_;
 wire clknet_1_0__leaf__04437_;
 wire clknet_1_0__leaf__04438_;
 wire clknet_1_0__leaf__04439_;
 wire clknet_1_0__leaf__04440_;
 wire clknet_1_0__leaf__04441_;
 wire clknet_1_0__leaf__04442_;
 wire clknet_1_0__leaf__04443_;
 wire clknet_1_0__leaf__04444_;
 wire clknet_1_0__leaf__04445_;
 wire clknet_1_0__leaf__04446_;
 wire clknet_1_0__leaf__04447_;
 wire clknet_1_0__leaf__04448_;
 wire clknet_1_0__leaf__04449_;
 wire clknet_1_0__leaf__04450_;
 wire clknet_1_0__leaf__04451_;
 wire clknet_1_0__leaf__04452_;
 wire clknet_1_0__leaf__04453_;
 wire clknet_1_0__leaf__04454_;
 wire clknet_1_0__leaf__04455_;
 wire clknet_1_0__leaf__04456_;
 wire clknet_1_0__leaf__04457_;
 wire clknet_1_0__leaf__04458_;
 wire clknet_1_0__leaf__04459_;
 wire clknet_1_0__leaf__04460_;
 wire clknet_1_0__leaf__04461_;
 wire clknet_1_0__leaf__04463_;
 wire clknet_1_0__leaf__04464_;
 wire clknet_1_0__leaf__04465_;
 wire clknet_1_0__leaf__04466_;
 wire clknet_1_0__leaf__04467_;
 wire clknet_1_0__leaf__04468_;
 wire clknet_1_0__leaf__04469_;
 wire clknet_1_0__leaf__04470_;
 wire clknet_1_0__leaf__04471_;
 wire clknet_1_0__leaf__04472_;
 wire clknet_1_0__leaf__04473_;
 wire clknet_1_0__leaf__04474_;
 wire clknet_1_0__leaf__04475_;
 wire clknet_1_0__leaf__04476_;
 wire clknet_1_0__leaf__04477_;
 wire clknet_1_0__leaf__04478_;
 wire clknet_1_0__leaf__04479_;
 wire clknet_1_0__leaf__04480_;
 wire clknet_1_0__leaf__04481_;
 wire clknet_1_0__leaf__04482_;
 wire clknet_1_0__leaf__04483_;
 wire clknet_1_0__leaf__04484_;
 wire clknet_1_0__leaf__04485_;
 wire clknet_1_0__leaf__04486_;
 wire clknet_1_0__leaf__04487_;
 wire clknet_1_0__leaf__04488_;
 wire clknet_1_0__leaf__04489_;
 wire clknet_1_0__leaf__04490_;
 wire clknet_1_0__leaf__04491_;
 wire clknet_1_0__leaf__04492_;
 wire clknet_1_0__leaf__04494_;
 wire clknet_1_0__leaf__04495_;
 wire clknet_1_0__leaf__04496_;
 wire clknet_1_0__leaf__04497_;
 wire clknet_1_0__leaf__04498_;
 wire clknet_1_0__leaf__04499_;
 wire clknet_1_0__leaf__04500_;
 wire clknet_1_0__leaf__04501_;
 wire clknet_1_0__leaf__04502_;
 wire clknet_1_0__leaf__04503_;
 wire clknet_1_0__leaf__04504_;
 wire clknet_1_0__leaf__04505_;
 wire clknet_1_0__leaf__04538_;
 wire clknet_1_0__leaf__04539_;
 wire clknet_1_0__leaf__04540_;
 wire clknet_1_0__leaf__04541_;
 wire clknet_1_0__leaf__04542_;
 wire clknet_1_0__leaf__04543_;
 wire clknet_1_0__leaf__04544_;
 wire clknet_1_0__leaf__04545_;
 wire clknet_1_0__leaf__04546_;
 wire clknet_1_0__leaf__04547_;
 wire clknet_1_0__leaf__04548_;
 wire clknet_1_0__leaf__04549_;
 wire clknet_1_0__leaf__04550_;
 wire clknet_1_0__leaf__04551_;
 wire clknet_1_0__leaf__04552_;
 wire clknet_1_0__leaf__04562_;
 wire clknet_1_0__leaf__04565_;
 wire clknet_1_0__leaf__04566_;
 wire clknet_1_0__leaf__04568_;
 wire clknet_1_0__leaf__04569_;
 wire clknet_1_0__leaf__04570_;
 wire clknet_1_0__leaf__04571_;
 wire clknet_1_0__leaf__04572_;
 wire clknet_1_0__leaf__04573_;
 wire clknet_1_0__leaf__04574_;
 wire clknet_1_0__leaf__04575_;
 wire clknet_1_0__leaf__04576_;
 wire clknet_1_0__leaf__04577_;
 wire clknet_1_0__leaf__04578_;
 wire clknet_1_0__leaf__04579_;
 wire clknet_1_0__leaf__04580_;
 wire clknet_1_0__leaf__04581_;
 wire clknet_1_0__leaf__04582_;
 wire clknet_1_0__leaf__04583_;
 wire clknet_1_0__leaf__04584_;
 wire clknet_1_0__leaf__04587_;
 wire clknet_1_0__leaf__04588_;
 wire clknet_1_0__leaf__04590_;
 wire clknet_1_0__leaf__04591_;
 wire clknet_1_0__leaf__04592_;
 wire clknet_1_0__leaf__04593_;
 wire clknet_1_0__leaf__04594_;
 wire clknet_1_0__leaf__04595_;
 wire clknet_1_0__leaf__04596_;
 wire clknet_1_0__leaf__04597_;
 wire clknet_1_0__leaf__04598_;
 wire clknet_1_0__leaf__04599_;
 wire clknet_1_0__leaf__04600_;
 wire clknet_1_0__leaf__04601_;
 wire clknet_1_0__leaf__04602_;
 wire clknet_1_0__leaf__04603_;
 wire clknet_1_0__leaf__04604_;
 wire clknet_1_0__leaf__04605_;
 wire clknet_1_0__leaf__04606_;
 wire clknet_1_0__leaf__04609_;
 wire clknet_1_0__leaf__04610_;
 wire clknet_1_0__leaf__04612_;
 wire clknet_1_0__leaf__04613_;
 wire clknet_1_0__leaf__04614_;
 wire clknet_1_0__leaf__04615_;
 wire clknet_1_0__leaf__04616_;
 wire clknet_1_0__leaf__04617_;
 wire clknet_1_0__leaf__04618_;
 wire clknet_1_0__leaf__04619_;
 wire clknet_1_0__leaf__04620_;
 wire clknet_1_0__leaf__04621_;
 wire clknet_1_0__leaf__04622_;
 wire clknet_1_0__leaf__04623_;
 wire clknet_1_0__leaf__04624_;
 wire clknet_1_0__leaf__04625_;
 wire clknet_1_0__leaf__04626_;
 wire clknet_1_0__leaf__04627_;
 wire clknet_1_0__leaf__04628_;
 wire clknet_1_0__leaf__04629_;
 wire clknet_1_0__leaf__04630_;
 wire clknet_1_0__leaf__04631_;
 wire clknet_1_0__leaf__04632_;
 wire clknet_1_0__leaf__04634_;
 wire clknet_1_0__leaf__04635_;
 wire clknet_1_0__leaf__04636_;
 wire clknet_1_0__leaf__04637_;
 wire clknet_1_0__leaf__04638_;
 wire clknet_1_0__leaf__04639_;
 wire clknet_1_0__leaf__04640_;
 wire clknet_1_0__leaf__04641_;
 wire clknet_1_0__leaf__04642_;
 wire clknet_1_0__leaf__04643_;
 wire clknet_1_0__leaf__04644_;
 wire clknet_1_0__leaf__04645_;
 wire clknet_1_0__leaf__04646_;
 wire clknet_1_0__leaf__04647_;
 wire clknet_1_0__leaf__04648_;
 wire clknet_1_0__leaf__04649_;
 wire clknet_1_0__leaf__04650_;
 wire clknet_1_0__leaf__04651_;
 wire clknet_1_0__leaf__04652_;
 wire clknet_1_0__leaf__04658_;
 wire clknet_1_0__leaf__04659_;
 wire clknet_1_0__leaf__04664_;
 wire clknet_1_0__leaf__04665_;
 wire clknet_1_0__leaf__04670_;
 wire clknet_1_0__leaf__04671_;
 wire clknet_1_0__leaf__04672_;
 wire clknet_1_0__leaf__04673_;
 wire clknet_1_0__leaf__04674_;
 wire clknet_1_0__leaf__04675_;
 wire clknet_1_0__leaf__04676_;
 wire clknet_1_0__leaf__04679_;
 wire clknet_1_0__leaf__04680_;
 wire clknet_1_0__leaf__04682_;
 wire clknet_1_0__leaf__04685_;
 wire clknet_1_0__leaf__04686_;
 wire clknet_1_0__leaf_user_clock1;
 wire clknet_1_0__leaf_user_clock2;
 wire clknet_1_1__leaf__04347_;
 wire clknet_1_1__leaf__04354_;
 wire clknet_1_1__leaf__04355_;
 wire clknet_1_1__leaf__04356_;
 wire clknet_1_1__leaf__04357_;
 wire clknet_1_1__leaf__04392_;
 wire clknet_1_1__leaf__04393_;
 wire clknet_1_1__leaf__04394_;
 wire clknet_1_1__leaf__04395_;
 wire clknet_1_1__leaf__04396_;
 wire clknet_1_1__leaf__04397_;
 wire clknet_1_1__leaf__04398_;
 wire clknet_1_1__leaf__04399_;
 wire clknet_1_1__leaf__04400_;
 wire clknet_1_1__leaf__04401_;
 wire clknet_1_1__leaf__04402_;
 wire clknet_1_1__leaf__04403_;
 wire clknet_1_1__leaf__04404_;
 wire clknet_1_1__leaf__04405_;
 wire clknet_1_1__leaf__04406_;
 wire clknet_1_1__leaf__04407_;
 wire clknet_1_1__leaf__04408_;
 wire clknet_1_1__leaf__04409_;
 wire clknet_1_1__leaf__04410_;
 wire clknet_1_1__leaf__04411_;
 wire clknet_1_1__leaf__04412_;
 wire clknet_1_1__leaf__04413_;
 wire clknet_1_1__leaf__04414_;
 wire clknet_1_1__leaf__04415_;
 wire clknet_1_1__leaf__04416_;
 wire clknet_1_1__leaf__04417_;
 wire clknet_1_1__leaf__04418_;
 wire clknet_1_1__leaf__04419_;
 wire clknet_1_1__leaf__04420_;
 wire clknet_1_1__leaf__04421_;
 wire clknet_1_1__leaf__04422_;
 wire clknet_1_1__leaf__04423_;
 wire clknet_1_1__leaf__04424_;
 wire clknet_1_1__leaf__04425_;
 wire clknet_1_1__leaf__04426_;
 wire clknet_1_1__leaf__04427_;
 wire clknet_1_1__leaf__04428_;
 wire clknet_1_1__leaf__04429_;
 wire clknet_1_1__leaf__04430_;
 wire clknet_1_1__leaf__04431_;
 wire clknet_1_1__leaf__04432_;
 wire clknet_1_1__leaf__04433_;
 wire clknet_1_1__leaf__04434_;
 wire clknet_1_1__leaf__04435_;
 wire clknet_1_1__leaf__04436_;
 wire clknet_1_1__leaf__04437_;
 wire clknet_1_1__leaf__04438_;
 wire clknet_1_1__leaf__04439_;
 wire clknet_1_1__leaf__04440_;
 wire clknet_1_1__leaf__04441_;
 wire clknet_1_1__leaf__04442_;
 wire clknet_1_1__leaf__04443_;
 wire clknet_1_1__leaf__04444_;
 wire clknet_1_1__leaf__04445_;
 wire clknet_1_1__leaf__04446_;
 wire clknet_1_1__leaf__04447_;
 wire clknet_1_1__leaf__04448_;
 wire clknet_1_1__leaf__04449_;
 wire clknet_1_1__leaf__04450_;
 wire clknet_1_1__leaf__04451_;
 wire clknet_1_1__leaf__04452_;
 wire clknet_1_1__leaf__04453_;
 wire clknet_1_1__leaf__04454_;
 wire clknet_1_1__leaf__04455_;
 wire clknet_1_1__leaf__04456_;
 wire clknet_1_1__leaf__04457_;
 wire clknet_1_1__leaf__04458_;
 wire clknet_1_1__leaf__04459_;
 wire clknet_1_1__leaf__04460_;
 wire clknet_1_1__leaf__04461_;
 wire clknet_1_1__leaf__04463_;
 wire clknet_1_1__leaf__04464_;
 wire clknet_1_1__leaf__04465_;
 wire clknet_1_1__leaf__04466_;
 wire clknet_1_1__leaf__04467_;
 wire clknet_1_1__leaf__04468_;
 wire clknet_1_1__leaf__04469_;
 wire clknet_1_1__leaf__04470_;
 wire clknet_1_1__leaf__04471_;
 wire clknet_1_1__leaf__04472_;
 wire clknet_1_1__leaf__04473_;
 wire clknet_1_1__leaf__04474_;
 wire clknet_1_1__leaf__04475_;
 wire clknet_1_1__leaf__04476_;
 wire clknet_1_1__leaf__04477_;
 wire clknet_1_1__leaf__04478_;
 wire clknet_1_1__leaf__04479_;
 wire clknet_1_1__leaf__04480_;
 wire clknet_1_1__leaf__04481_;
 wire clknet_1_1__leaf__04482_;
 wire clknet_1_1__leaf__04483_;
 wire clknet_1_1__leaf__04484_;
 wire clknet_1_1__leaf__04485_;
 wire clknet_1_1__leaf__04486_;
 wire clknet_1_1__leaf__04487_;
 wire clknet_1_1__leaf__04488_;
 wire clknet_1_1__leaf__04489_;
 wire clknet_1_1__leaf__04490_;
 wire clknet_1_1__leaf__04491_;
 wire clknet_1_1__leaf__04492_;
 wire clknet_1_1__leaf__04494_;
 wire clknet_1_1__leaf__04495_;
 wire clknet_1_1__leaf__04496_;
 wire clknet_1_1__leaf__04497_;
 wire clknet_1_1__leaf__04498_;
 wire clknet_1_1__leaf__04499_;
 wire clknet_1_1__leaf__04500_;
 wire clknet_1_1__leaf__04501_;
 wire clknet_1_1__leaf__04502_;
 wire clknet_1_1__leaf__04503_;
 wire clknet_1_1__leaf__04504_;
 wire clknet_1_1__leaf__04505_;
 wire clknet_1_1__leaf__04538_;
 wire clknet_1_1__leaf__04539_;
 wire clknet_1_1__leaf__04540_;
 wire clknet_1_1__leaf__04541_;
 wire clknet_1_1__leaf__04542_;
 wire clknet_1_1__leaf__04543_;
 wire clknet_1_1__leaf__04544_;
 wire clknet_1_1__leaf__04545_;
 wire clknet_1_1__leaf__04546_;
 wire clknet_1_1__leaf__04547_;
 wire clknet_1_1__leaf__04548_;
 wire clknet_1_1__leaf__04549_;
 wire clknet_1_1__leaf__04550_;
 wire clknet_1_1__leaf__04551_;
 wire clknet_1_1__leaf__04552_;
 wire clknet_1_1__leaf__04562_;
 wire clknet_1_1__leaf__04565_;
 wire clknet_1_1__leaf__04566_;
 wire clknet_1_1__leaf__04568_;
 wire clknet_1_1__leaf__04569_;
 wire clknet_1_1__leaf__04570_;
 wire clknet_1_1__leaf__04571_;
 wire clknet_1_1__leaf__04572_;
 wire clknet_1_1__leaf__04573_;
 wire clknet_1_1__leaf__04574_;
 wire clknet_1_1__leaf__04575_;
 wire clknet_1_1__leaf__04576_;
 wire clknet_1_1__leaf__04577_;
 wire clknet_1_1__leaf__04578_;
 wire clknet_1_1__leaf__04579_;
 wire clknet_1_1__leaf__04580_;
 wire clknet_1_1__leaf__04581_;
 wire clknet_1_1__leaf__04582_;
 wire clknet_1_1__leaf__04583_;
 wire clknet_1_1__leaf__04584_;
 wire clknet_1_1__leaf__04587_;
 wire clknet_1_1__leaf__04588_;
 wire clknet_1_1__leaf__04590_;
 wire clknet_1_1__leaf__04591_;
 wire clknet_1_1__leaf__04592_;
 wire clknet_1_1__leaf__04593_;
 wire clknet_1_1__leaf__04594_;
 wire clknet_1_1__leaf__04595_;
 wire clknet_1_1__leaf__04596_;
 wire clknet_1_1__leaf__04597_;
 wire clknet_1_1__leaf__04598_;
 wire clknet_1_1__leaf__04599_;
 wire clknet_1_1__leaf__04600_;
 wire clknet_1_1__leaf__04601_;
 wire clknet_1_1__leaf__04602_;
 wire clknet_1_1__leaf__04603_;
 wire clknet_1_1__leaf__04604_;
 wire clknet_1_1__leaf__04605_;
 wire clknet_1_1__leaf__04606_;
 wire clknet_1_1__leaf__04609_;
 wire clknet_1_1__leaf__04610_;
 wire clknet_1_1__leaf__04612_;
 wire clknet_1_1__leaf__04613_;
 wire clknet_1_1__leaf__04614_;
 wire clknet_1_1__leaf__04615_;
 wire clknet_1_1__leaf__04616_;
 wire clknet_1_1__leaf__04617_;
 wire clknet_1_1__leaf__04618_;
 wire clknet_1_1__leaf__04619_;
 wire clknet_1_1__leaf__04620_;
 wire clknet_1_1__leaf__04621_;
 wire clknet_1_1__leaf__04622_;
 wire clknet_1_1__leaf__04623_;
 wire clknet_1_1__leaf__04624_;
 wire clknet_1_1__leaf__04625_;
 wire clknet_1_1__leaf__04626_;
 wire clknet_1_1__leaf__04627_;
 wire clknet_1_1__leaf__04628_;
 wire clknet_1_1__leaf__04629_;
 wire clknet_1_1__leaf__04630_;
 wire clknet_1_1__leaf__04631_;
 wire clknet_1_1__leaf__04632_;
 wire clknet_1_1__leaf__04634_;
 wire clknet_1_1__leaf__04635_;
 wire clknet_1_1__leaf__04636_;
 wire clknet_1_1__leaf__04637_;
 wire clknet_1_1__leaf__04638_;
 wire clknet_1_1__leaf__04639_;
 wire clknet_1_1__leaf__04640_;
 wire clknet_1_1__leaf__04641_;
 wire clknet_1_1__leaf__04642_;
 wire clknet_1_1__leaf__04643_;
 wire clknet_1_1__leaf__04644_;
 wire clknet_1_1__leaf__04645_;
 wire clknet_1_1__leaf__04646_;
 wire clknet_1_1__leaf__04647_;
 wire clknet_1_1__leaf__04648_;
 wire clknet_1_1__leaf__04649_;
 wire clknet_1_1__leaf__04650_;
 wire clknet_1_1__leaf__04651_;
 wire clknet_1_1__leaf__04652_;
 wire clknet_1_1__leaf__04658_;
 wire clknet_1_1__leaf__04659_;
 wire clknet_1_1__leaf__04664_;
 wire clknet_1_1__leaf__04665_;
 wire clknet_1_1__leaf__04670_;
 wire clknet_1_1__leaf__04671_;
 wire clknet_1_1__leaf__04672_;
 wire clknet_1_1__leaf__04673_;
 wire clknet_1_1__leaf__04674_;
 wire clknet_1_1__leaf__04675_;
 wire clknet_1_1__leaf__04676_;
 wire clknet_1_1__leaf__04679_;
 wire clknet_1_1__leaf__04680_;
 wire clknet_1_1__leaf__04682_;
 wire clknet_1_1__leaf__04685_;
 wire clknet_1_1__leaf__04686_;
 wire clknet_1_1__leaf_user_clock1;
 wire clknet_1_1__leaf_user_clock2;
 wire clknet_2_0_0_mclk;
 wire clknet_2_0__leaf__04353_;
 wire clknet_2_0__leaf__04358_;
 wire clknet_2_0__leaf__04359_;
 wire clknet_2_0__leaf__04493_;
 wire clknet_2_0__leaf__04564_;
 wire clknet_2_0__leaf__04567_;
 wire clknet_2_0__leaf__04586_;
 wire clknet_2_0__leaf__04589_;
 wire clknet_2_0__leaf__04608_;
 wire clknet_2_0__leaf__04611_;
 wire clknet_2_0__leaf__04633_;
 wire clknet_2_0__leaf__04653_;
 wire clknet_2_1_0_mclk;
 wire clknet_2_1__leaf__04353_;
 wire clknet_2_1__leaf__04358_;
 wire clknet_2_1__leaf__04359_;
 wire clknet_2_1__leaf__04493_;
 wire clknet_2_1__leaf__04564_;
 wire clknet_2_1__leaf__04567_;
 wire clknet_2_1__leaf__04586_;
 wire clknet_2_1__leaf__04589_;
 wire clknet_2_1__leaf__04608_;
 wire clknet_2_1__leaf__04611_;
 wire clknet_2_1__leaf__04633_;
 wire clknet_2_1__leaf__04653_;
 wire clknet_2_2_0_mclk;
 wire clknet_2_2__leaf__04353_;
 wire clknet_2_2__leaf__04358_;
 wire clknet_2_2__leaf__04359_;
 wire clknet_2_2__leaf__04493_;
 wire clknet_2_2__leaf__04564_;
 wire clknet_2_2__leaf__04567_;
 wire clknet_2_2__leaf__04586_;
 wire clknet_2_2__leaf__04589_;
 wire clknet_2_2__leaf__04608_;
 wire clknet_2_2__leaf__04611_;
 wire clknet_2_2__leaf__04633_;
 wire clknet_2_2__leaf__04653_;
 wire clknet_2_3_0_mclk;
 wire clknet_2_3__leaf__04353_;
 wire clknet_2_3__leaf__04358_;
 wire clknet_2_3__leaf__04359_;
 wire clknet_2_3__leaf__04493_;
 wire clknet_2_3__leaf__04564_;
 wire clknet_2_3__leaf__04567_;
 wire clknet_2_3__leaf__04586_;
 wire clknet_2_3__leaf__04589_;
 wire clknet_2_3__leaf__04608_;
 wire clknet_2_3__leaf__04611_;
 wire clknet_2_3__leaf__04633_;
 wire clknet_2_3__leaf__04653_;
 wire clknet_4_0__leaf_mclk;
 wire clknet_4_10__leaf_mclk;
 wire clknet_4_11__leaf_mclk;
 wire clknet_4_12__leaf_mclk;
 wire clknet_4_13__leaf_mclk;
 wire clknet_4_14__leaf_mclk;
 wire clknet_4_15__leaf_mclk;
 wire clknet_4_1__leaf_mclk;
 wire clknet_4_2__leaf_mclk;
 wire clknet_4_3__leaf_mclk;
 wire clknet_4_4__leaf_mclk;
 wire clknet_4_5__leaf_mclk;
 wire clknet_4_6__leaf_mclk;
 wire clknet_4_7__leaf_mclk;
 wire clknet_4_8__leaf_mclk;
 wire clknet_4_9__leaf_mclk;
 wire clknet_leaf_0_mclk;
 wire clknet_leaf_100_mclk;
 wire clknet_leaf_102_mclk;
 wire clknet_leaf_103_mclk;
 wire clknet_leaf_104_mclk;
 wire clknet_leaf_105_mclk;
 wire clknet_leaf_106_mclk;
 wire clknet_leaf_107_mclk;
 wire clknet_leaf_109_mclk;
 wire clknet_leaf_10_mclk;
 wire clknet_leaf_110_mclk;
 wire clknet_leaf_111_mclk;
 wire clknet_leaf_112_mclk;
 wire clknet_leaf_113_mclk;
 wire clknet_leaf_114_mclk;
 wire clknet_leaf_115_mclk;
 wire clknet_leaf_116_mclk;
 wire clknet_leaf_117_mclk;
 wire clknet_leaf_118_mclk;
 wire clknet_leaf_11_mclk;
 wire clknet_leaf_120_mclk;
 wire clknet_leaf_122_mclk;
 wire clknet_leaf_123_mclk;
 wire clknet_leaf_124_mclk;
 wire clknet_leaf_126_mclk;
 wire clknet_leaf_127_mclk;
 wire clknet_leaf_128_mclk;
 wire clknet_leaf_12_mclk;
 wire clknet_leaf_13_mclk;
 wire clknet_leaf_14_mclk;
 wire clknet_leaf_15_mclk;
 wire clknet_leaf_16_mclk;
 wire clknet_leaf_17_mclk;
 wire clknet_leaf_19_mclk;
 wire clknet_leaf_1_mclk;
 wire clknet_leaf_20_mclk;
 wire clknet_leaf_21_mclk;
 wire clknet_leaf_22_mclk;
 wire clknet_leaf_23_mclk;
 wire clknet_leaf_24_mclk;
 wire clknet_leaf_25_mclk;
 wire clknet_leaf_26_mclk;
 wire clknet_leaf_28_mclk;
 wire clknet_leaf_29_mclk;
 wire clknet_leaf_2_mclk;
 wire clknet_leaf_30_mclk;
 wire clknet_leaf_31_mclk;
 wire clknet_leaf_32_mclk;
 wire clknet_leaf_33_mclk;
 wire clknet_leaf_34_mclk;
 wire clknet_leaf_35_mclk;
 wire clknet_leaf_36_mclk;
 wire clknet_leaf_37_mclk;
 wire clknet_leaf_38_mclk;
 wire clknet_leaf_39_mclk;
 wire clknet_leaf_40_mclk;
 wire clknet_leaf_41_mclk;
 wire clknet_leaf_42_mclk;
 wire clknet_leaf_43_mclk;
 wire clknet_leaf_44_mclk;
 wire clknet_leaf_45_mclk;
 wire clknet_leaf_46_mclk;
 wire clknet_leaf_47_mclk;
 wire clknet_leaf_48_mclk;
 wire clknet_leaf_4_mclk;
 wire clknet_leaf_51_mclk;
 wire clknet_leaf_53_mclk;
 wire clknet_leaf_54_mclk;
 wire clknet_leaf_55_mclk;
 wire clknet_leaf_56_mclk;
 wire clknet_leaf_58_mclk;
 wire clknet_leaf_5_mclk;
 wire clknet_leaf_60_mclk;
 wire clknet_leaf_62_mclk;
 wire clknet_leaf_63_mclk;
 wire clknet_leaf_65_mclk;
 wire clknet_leaf_66_mclk;
 wire clknet_leaf_67_mclk;
 wire clknet_leaf_69_mclk;
 wire clknet_leaf_6_mclk;
 wire clknet_leaf_70_mclk;
 wire clknet_leaf_72_mclk;
 wire clknet_leaf_73_mclk;
 wire clknet_leaf_74_mclk;
 wire clknet_leaf_75_mclk;
 wire clknet_leaf_76_mclk;
 wire clknet_leaf_77_mclk;
 wire clknet_leaf_78_mclk;
 wire clknet_leaf_79_mclk;
 wire clknet_leaf_7_mclk;
 wire clknet_leaf_80_mclk;
 wire clknet_leaf_81_mclk;
 wire clknet_leaf_82_mclk;
 wire clknet_leaf_83_mclk;
 wire clknet_leaf_84_mclk;
 wire clknet_leaf_85_mclk;
 wire clknet_leaf_86_mclk;
 wire clknet_leaf_87_mclk;
 wire clknet_leaf_88_mclk;
 wire clknet_leaf_89_mclk;
 wire clknet_leaf_8_mclk;
 wire clknet_leaf_90_mclk;
 wire clknet_leaf_91_mclk;
 wire clknet_leaf_92_mclk;
 wire clknet_leaf_93_mclk;
 wire clknet_leaf_94_mclk;
 wire clknet_leaf_95_mclk;
 wire clknet_leaf_96_mclk;
 wire clknet_leaf_97_mclk;
 wire clknet_leaf_99_mclk;
 wire clknet_leaf_9_mclk;
 wire net1;
 wire net10;
 wire net100;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net101;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net102;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net103;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net104;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net105;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net106;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net107;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net108;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net109;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net11;
 wire net110;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net111;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net112;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net113;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net114;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net115;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net116;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net117;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net118;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net119;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;
 wire net1198;
 wire net1199;
 wire net12;
 wire net120;
 wire net1200;
 wire net1201;
 wire net1202;
 wire net1203;
 wire net1204;
 wire net1205;
 wire net1206;
 wire net1207;
 wire net1208;
 wire net1209;
 wire net121;
 wire net1210;
 wire net1211;
 wire net1212;
 wire net1213;
 wire net1214;
 wire net1215;
 wire net1216;
 wire net1217;
 wire net1218;
 wire net1219;
 wire net122;
 wire net1220;
 wire net1221;
 wire net1222;
 wire net1223;
 wire net1224;
 wire net1225;
 wire net1226;
 wire net1227;
 wire net1228;
 wire net1229;
 wire net123;
 wire net1230;
 wire net1231;
 wire net1232;
 wire net1233;
 wire net1234;
 wire net1235;
 wire net1236;
 wire net1237;
 wire net1238;
 wire net1239;
 wire net124;
 wire net1240;
 wire net1241;
 wire net1242;
 wire net1243;
 wire net1244;
 wire net1245;
 wire net1246;
 wire net1247;
 wire net1248;
 wire net1249;
 wire net125;
 wire net1250;
 wire net1251;
 wire net1252;
 wire net1253;
 wire net1254;
 wire net1255;
 wire net1256;
 wire net1257;
 wire net1258;
 wire net1259;
 wire net126;
 wire net1260;
 wire net1261;
 wire net1262;
 wire net1263;
 wire net1264;
 wire net1265;
 wire net1266;
 wire net1267;
 wire net1268;
 wire net1269;
 wire net127;
 wire net1270;
 wire net1271;
 wire net1272;
 wire net1273;
 wire net1274;
 wire net1275;
 wire net1276;
 wire net1277;
 wire net1278;
 wire net1279;
 wire net128;
 wire net1280;
 wire net1281;
 wire net1282;
 wire net1283;
 wire net1284;
 wire net1285;
 wire net1286;
 wire net1287;
 wire net1288;
 wire net1289;
 wire net129;
 wire net1290;
 wire net1291;
 wire net1292;
 wire net1293;
 wire net1294;
 wire net1295;
 wire net1296;
 wire net1297;
 wire net1298;
 wire net1299;
 wire net13;
 wire net130;
 wire net1300;
 wire net1301;
 wire net1302;
 wire net1303;
 wire net1304;
 wire net1305;
 wire net1306;
 wire net1307;
 wire net1308;
 wire net1309;
 wire net131;
 wire net1310;
 wire net1311;
 wire net1312;
 wire net1313;
 wire net1314;
 wire net1315;
 wire net1316;
 wire net1317;
 wire net1318;
 wire net1319;
 wire net132;
 wire net1320;
 wire net1321;
 wire net1322;
 wire net1323;
 wire net1324;
 wire net1325;
 wire net1326;
 wire net1327;
 wire net1328;
 wire net1329;
 wire net133;
 wire net1330;
 wire net1331;
 wire net1332;
 wire net1333;
 wire net1334;
 wire net1335;
 wire net1336;
 wire net1337;
 wire net1338;
 wire net1339;
 wire net134;
 wire net1340;
 wire net1341;
 wire net1342;
 wire net1343;
 wire net1344;
 wire net1345;
 wire net1346;
 wire net1347;
 wire net1348;
 wire net1349;
 wire net135;
 wire net1350;
 wire net1351;
 wire net1352;
 wire net1353;
 wire net1354;
 wire net1355;
 wire net1356;
 wire net1357;
 wire net1358;
 wire net1359;
 wire net136;
 wire net1360;
 wire net1361;
 wire net1362;
 wire net1363;
 wire net1364;
 wire net1365;
 wire net1366;
 wire net1367;
 wire net1368;
 wire net1369;
 wire net137;
 wire net1370;
 wire net1371;
 wire net1372;
 wire net1373;
 wire net1374;
 wire net1375;
 wire net1376;
 wire net1377;
 wire net1378;
 wire net1379;
 wire net138;
 wire net1380;
 wire net1381;
 wire net1382;
 wire net1383;
 wire net1384;
 wire net1385;
 wire net1386;
 wire net1387;
 wire net1388;
 wire net1389;
 wire net139;
 wire net1390;
 wire net1391;
 wire net1392;
 wire net1393;
 wire net1394;
 wire net1395;
 wire net1396;
 wire net1397;
 wire net1398;
 wire net1399;
 wire net14;
 wire net140;
 wire net1400;
 wire net1401;
 wire net1402;
 wire net1403;
 wire net1404;
 wire net1405;
 wire net1406;
 wire net1407;
 wire net1408;
 wire net1409;
 wire net141;
 wire net1410;
 wire net1411;
 wire net1412;
 wire net1413;
 wire net1414;
 wire net1415;
 wire net1416;
 wire net1417;
 wire net1418;
 wire net1419;
 wire net142;
 wire net1420;
 wire net1421;
 wire net1422;
 wire net1423;
 wire net1424;
 wire net1425;
 wire net1426;
 wire net1427;
 wire net1428;
 wire net1429;
 wire net143;
 wire net1430;
 wire net1431;
 wire net1432;
 wire net1433;
 wire net1434;
 wire net1435;
 wire net1436;
 wire net1437;
 wire net1438;
 wire net1439;
 wire net144;
 wire net1440;
 wire net1441;
 wire net1442;
 wire net1443;
 wire net1444;
 wire net1445;
 wire net1446;
 wire net1447;
 wire net1448;
 wire net1449;
 wire net145;
 wire net1450;
 wire net1451;
 wire net1452;
 wire net1453;
 wire net1454;
 wire net1455;
 wire net1456;
 wire net1457;
 wire net1458;
 wire net1459;
 wire net146;
 wire net1460;
 wire net1461;
 wire net1462;
 wire net1463;
 wire net1464;
 wire net1465;
 wire net1466;
 wire net1467;
 wire net1468;
 wire net1469;
 wire net147;
 wire net1470;
 wire net1471;
 wire net1472;
 wire net1473;
 wire net1474;
 wire net1475;
 wire net1476;
 wire net1477;
 wire net1478;
 wire net1479;
 wire net148;
 wire net1480;
 wire net1481;
 wire net1482;
 wire net1483;
 wire net1484;
 wire net1485;
 wire net1486;
 wire net1487;
 wire net1488;
 wire net1489;
 wire net149;
 wire net1490;
 wire net1491;
 wire net1492;
 wire net1493;
 wire net1494;
 wire net1495;
 wire net1496;
 wire net1497;
 wire net1498;
 wire net1499;
 wire net15;
 wire net150;
 wire net1500;
 wire net1501;
 wire net1502;
 wire net1503;
 wire net1504;
 wire net1505;
 wire net1506;
 wire net1507;
 wire net1508;
 wire net1509;
 wire net151;
 wire net1510;
 wire net1511;
 wire net1512;
 wire net1513;
 wire net1514;
 wire net1515;
 wire net1516;
 wire net1517;
 wire net1518;
 wire net1519;
 wire net152;
 wire net1520;
 wire net1521;
 wire net1522;
 wire net1523;
 wire net1524;
 wire net1525;
 wire net1526;
 wire net1527;
 wire net1528;
 wire net1529;
 wire net153;
 wire net1530;
 wire net1531;
 wire net1532;
 wire net1533;
 wire net1534;
 wire net1535;
 wire net1536;
 wire net1537;
 wire net1538;
 wire net1539;
 wire net154;
 wire net1540;
 wire net1541;
 wire net1542;
 wire net1543;
 wire net1544;
 wire net1545;
 wire net1546;
 wire net1547;
 wire net1548;
 wire net1549;
 wire net155;
 wire net1550;
 wire net1551;
 wire net1552;
 wire net1553;
 wire net1554;
 wire net1555;
 wire net1556;
 wire net1557;
 wire net1558;
 wire net1559;
 wire net156;
 wire net1560;
 wire net1561;
 wire net1562;
 wire net1563;
 wire net1564;
 wire net1565;
 wire net1566;
 wire net1567;
 wire net1568;
 wire net1569;
 wire net157;
 wire net1570;
 wire net1571;
 wire net1572;
 wire net1573;
 wire net1574;
 wire net1575;
 wire net1576;
 wire net1577;
 wire net1578;
 wire net1579;
 wire net158;
 wire net1580;
 wire net1581;
 wire net1582;
 wire net1583;
 wire net1584;
 wire net1585;
 wire net1586;
 wire net1587;
 wire net1588;
 wire net1589;
 wire net159;
 wire net1590;
 wire net1591;
 wire net1592;
 wire net1593;
 wire net1594;
 wire net1595;
 wire net1596;
 wire net1597;
 wire net1598;
 wire net1599;
 wire net16;
 wire net160;
 wire net1600;
 wire net1601;
 wire net1602;
 wire net1603;
 wire net1604;
 wire net1605;
 wire net1606;
 wire net1607;
 wire net1608;
 wire net1609;
 wire net161;
 wire net1610;
 wire net1611;
 wire net1612;
 wire net1613;
 wire net1614;
 wire net1615;
 wire net1616;
 wire net1617;
 wire net1618;
 wire net1619;
 wire net162;
 wire net1620;
 wire net1621;
 wire net1622;
 wire net1623;
 wire net1624;
 wire net1625;
 wire net1626;
 wire net1627;
 wire net1628;
 wire net1629;
 wire net163;
 wire net1630;
 wire net1631;
 wire net1632;
 wire net1633;
 wire net1634;
 wire net1635;
 wire net1636;
 wire net1637;
 wire net1638;
 wire net1639;
 wire net164;
 wire net1640;
 wire net1641;
 wire net1642;
 wire net1643;
 wire net1644;
 wire net1645;
 wire net1646;
 wire net1647;
 wire net1648;
 wire net1649;
 wire net165;
 wire net1650;
 wire net1651;
 wire net1652;
 wire net1653;
 wire net1654;
 wire net1655;
 wire net1656;
 wire net166;
 wire net167;
 wire net168;
 wire net1689;
 wire net169;
 wire net1690;
 wire net1691;
 wire net1692;
 wire net1693;
 wire net1694;
 wire net1695;
 wire net1696;
 wire net1697;
 wire net1698;
 wire net1699;
 wire net17;
 wire net170;
 wire net1700;
 wire net1701;
 wire net1702;
 wire net1703;
 wire net1704;
 wire net1705;
 wire net1706;
 wire net1707;
 wire net1708;
 wire net1709;
 wire net171;
 wire net1710;
 wire net1711;
 wire net1712;
 wire net1713;
 wire net1714;
 wire net1715;
 wire net1716;
 wire net1717;
 wire net1718;
 wire net1719;
 wire net172;
 wire net1720;
 wire net1721;
 wire net1722;
 wire net1723;
 wire net1724;
 wire net1725;
 wire net1726;
 wire net1727;
 wire net1728;
 wire net1729;
 wire net173;
 wire net1730;
 wire net1731;
 wire net1732;
 wire net1733;
 wire net1734;
 wire net1735;
 wire net1736;
 wire net1737;
 wire net1738;
 wire net1739;
 wire net174;
 wire net1740;
 wire net1741;
 wire net1742;
 wire net1743;
 wire net1744;
 wire net1745;
 wire net1746;
 wire net1747;
 wire net1748;
 wire net1749;
 wire net175;
 wire net1750;
 wire net1751;
 wire net1752;
 wire net1753;
 wire net1754;
 wire net1755;
 wire net1756;
 wire net1757;
 wire net1758;
 wire net1759;
 wire net176;
 wire net1760;
 wire net1761;
 wire net1762;
 wire net1763;
 wire net1764;
 wire net1765;
 wire net1766;
 wire net1767;
 wire net1768;
 wire net1769;
 wire net177;
 wire net1770;
 wire net1771;
 wire net1772;
 wire net1773;
 wire net1774;
 wire net1775;
 wire net1776;
 wire net1777;
 wire net1778;
 wire net1779;
 wire net178;
 wire net1780;
 wire net1781;
 wire net1782;
 wire net1783;
 wire net1784;
 wire net1785;
 wire net1786;
 wire net1787;
 wire net1788;
 wire net1789;
 wire net179;
 wire net1790;
 wire net1791;
 wire net1792;
 wire net1793;
 wire net1794;
 wire net1795;
 wire net1796;
 wire net1797;
 wire net1798;
 wire net1799;
 wire net18;
 wire net180;
 wire net1800;
 wire net1801;
 wire net1802;
 wire net1803;
 wire net1804;
 wire net1805;
 wire net1806;
 wire net1807;
 wire net1808;
 wire net1809;
 wire net181;
 wire net1810;
 wire net1811;
 wire net1812;
 wire net1813;
 wire net1814;
 wire net1815;
 wire net1816;
 wire net1817;
 wire net1818;
 wire net1819;
 wire net182;
 wire net1820;
 wire net1821;
 wire net1822;
 wire net1823;
 wire net1824;
 wire net1825;
 wire net1826;
 wire net1827;
 wire net1828;
 wire net1829;
 wire net183;
 wire net1830;
 wire net1831;
 wire net1832;
 wire net1833;
 wire net1834;
 wire net1835;
 wire net1836;
 wire net1837;
 wire net1838;
 wire net1839;
 wire net184;
 wire net1840;
 wire net1841;
 wire net1842;
 wire net1843;
 wire net1844;
 wire net1845;
 wire net1846;
 wire net1847;
 wire net1848;
 wire net1849;
 wire net185;
 wire net1850;
 wire net1851;
 wire net1852;
 wire net1853;
 wire net1854;
 wire net1855;
 wire net1856;
 wire net1857;
 wire net1858;
 wire net1859;
 wire net186;
 wire net1860;
 wire net1861;
 wire net1862;
 wire net1863;
 wire net1864;
 wire net1865;
 wire net1866;
 wire net1867;
 wire net1868;
 wire net1869;
 wire net187;
 wire net1870;
 wire net1871;
 wire net1872;
 wire net1873;
 wire net1874;
 wire net1875;
 wire net1876;
 wire net1877;
 wire net1878;
 wire net1879;
 wire net188;
 wire net1880;
 wire net1881;
 wire net1882;
 wire net1883;
 wire net1884;
 wire net1885;
 wire net1886;
 wire net1887;
 wire net1888;
 wire net1889;
 wire net189;
 wire net1890;
 wire net1891;
 wire net1892;
 wire net1893;
 wire net1894;
 wire net1895;
 wire net1896;
 wire net1897;
 wire net1898;
 wire net1899;
 wire net19;
 wire net190;
 wire net1900;
 wire net1901;
 wire net1902;
 wire net1903;
 wire net1904;
 wire net1905;
 wire net1906;
 wire net1907;
 wire net1908;
 wire net1909;
 wire net191;
 wire net1910;
 wire net1911;
 wire net1912;
 wire net1913;
 wire net1914;
 wire net1915;
 wire net1916;
 wire net1917;
 wire net1918;
 wire net1919;
 wire net192;
 wire net1920;
 wire net1921;
 wire net1922;
 wire net1923;
 wire net1924;
 wire net1925;
 wire net1926;
 wire net1927;
 wire net1928;
 wire net1929;
 wire net193;
 wire net1930;
 wire net1931;
 wire net1932;
 wire net1933;
 wire net1934;
 wire net1935;
 wire net1936;
 wire net1937;
 wire net1938;
 wire net1939;
 wire net194;
 wire net1940;
 wire net1941;
 wire net1942;
 wire net1943;
 wire net1944;
 wire net1945;
 wire net1946;
 wire net1947;
 wire net1948;
 wire net1949;
 wire net195;
 wire net1950;
 wire net1951;
 wire net1952;
 wire net1953;
 wire net1954;
 wire net1955;
 wire net1956;
 wire net1957;
 wire net1958;
 wire net1959;
 wire net196;
 wire net1960;
 wire net1961;
 wire net1962;
 wire net1963;
 wire net1964;
 wire net1965;
 wire net1966;
 wire net1967;
 wire net1968;
 wire net1969;
 wire net197;
 wire net1970;
 wire net1971;
 wire net1972;
 wire net1973;
 wire net1974;
 wire net1975;
 wire net1976;
 wire net1977;
 wire net1978;
 wire net1979;
 wire net198;
 wire net1980;
 wire net1981;
 wire net1982;
 wire net1983;
 wire net1984;
 wire net1985;
 wire net1986;
 wire net1987;
 wire net1988;
 wire net1989;
 wire net199;
 wire net1990;
 wire net1991;
 wire net1992;
 wire net1993;
 wire net1994;
 wire net1995;
 wire net1996;
 wire net1997;
 wire net1998;
 wire net1999;
 wire net2;
 wire net20;
 wire net200;
 wire net2000;
 wire net2001;
 wire net2002;
 wire net2003;
 wire net2004;
 wire net2005;
 wire net2006;
 wire net2007;
 wire net2008;
 wire net2009;
 wire net201;
 wire net2010;
 wire net2011;
 wire net2012;
 wire net2013;
 wire net2014;
 wire net2015;
 wire net2016;
 wire net2017;
 wire net2018;
 wire net2019;
 wire net202;
 wire net2020;
 wire net2021;
 wire net2022;
 wire net2023;
 wire net2024;
 wire net2025;
 wire net2026;
 wire net2027;
 wire net2028;
 wire net2029;
 wire net203;
 wire net2030;
 wire net2031;
 wire net2032;
 wire net2033;
 wire net2034;
 wire net2035;
 wire net2036;
 wire net2037;
 wire net2038;
 wire net2039;
 wire net204;
 wire net2040;
 wire net2041;
 wire net2042;
 wire net2043;
 wire net2044;
 wire net2045;
 wire net2046;
 wire net2047;
 wire net2048;
 wire net2049;
 wire net205;
 wire net2050;
 wire net2051;
 wire net2052;
 wire net2053;
 wire net2054;
 wire net2055;
 wire net2056;
 wire net2057;
 wire net2058;
 wire net2059;
 wire net206;
 wire net2060;
 wire net2061;
 wire net2062;
 wire net2063;
 wire net2064;
 wire net2065;
 wire net2066;
 wire net2067;
 wire net2068;
 wire net2069;
 wire net207;
 wire net2070;
 wire net2071;
 wire net2072;
 wire net2073;
 wire net2074;
 wire net2075;
 wire net2076;
 wire net2077;
 wire net2078;
 wire net2079;
 wire net208;
 wire net2080;
 wire net2081;
 wire net2082;
 wire net2083;
 wire net2084;
 wire net2085;
 wire net2086;
 wire net2087;
 wire net2088;
 wire net2089;
 wire net209;
 wire net2090;
 wire net2091;
 wire net2092;
 wire net2093;
 wire net2094;
 wire net2095;
 wire net2096;
 wire net2097;
 wire net2098;
 wire net2099;
 wire net21;
 wire net210;
 wire net2100;
 wire net2101;
 wire net2102;
 wire net2103;
 wire net2104;
 wire net2105;
 wire net2106;
 wire net2107;
 wire net2108;
 wire net2109;
 wire net211;
 wire net2110;
 wire net2111;
 wire net2112;
 wire net2113;
 wire net2114;
 wire net2115;
 wire net2116;
 wire net2117;
 wire net2118;
 wire net2119;
 wire net212;
 wire net2120;
 wire net2121;
 wire net2122;
 wire net2123;
 wire net2124;
 wire net2125;
 wire net2126;
 wire net2127;
 wire net2128;
 wire net2129;
 wire net213;
 wire net2130;
 wire net2131;
 wire net2132;
 wire net2133;
 wire net2134;
 wire net2135;
 wire net2136;
 wire net2137;
 wire net2138;
 wire net2139;
 wire net214;
 wire net2140;
 wire net2141;
 wire net2142;
 wire net2143;
 wire net2144;
 wire net2145;
 wire net2146;
 wire net2147;
 wire net2148;
 wire net2149;
 wire net215;
 wire net2150;
 wire net2151;
 wire net2152;
 wire net2153;
 wire net2154;
 wire net2155;
 wire net2156;
 wire net2157;
 wire net2158;
 wire net2159;
 wire net216;
 wire net2160;
 wire net2161;
 wire net2162;
 wire net2163;
 wire net2164;
 wire net2165;
 wire net2166;
 wire net2167;
 wire net2168;
 wire net2169;
 wire net217;
 wire net2170;
 wire net2171;
 wire net2172;
 wire net2173;
 wire net2174;
 wire net2175;
 wire net2176;
 wire net2177;
 wire net2178;
 wire net2179;
 wire net218;
 wire net2180;
 wire net2181;
 wire net2182;
 wire net2183;
 wire net2184;
 wire net2185;
 wire net2186;
 wire net2187;
 wire net2188;
 wire net2189;
 wire net219;
 wire net2190;
 wire net2191;
 wire net2192;
 wire net2193;
 wire net2194;
 wire net2195;
 wire net2196;
 wire net2197;
 wire net2198;
 wire net2199;
 wire net22;
 wire net220;
 wire net2200;
 wire net2201;
 wire net2202;
 wire net2203;
 wire net2204;
 wire net2205;
 wire net2206;
 wire net2207;
 wire net2208;
 wire net2209;
 wire net221;
 wire net2210;
 wire net2211;
 wire net2212;
 wire net2213;
 wire net2214;
 wire net2215;
 wire net2216;
 wire net2217;
 wire net2218;
 wire net2219;
 wire net222;
 wire net2220;
 wire net2221;
 wire net2222;
 wire net2223;
 wire net2224;
 wire net2225;
 wire net2226;
 wire net2227;
 wire net2228;
 wire net2229;
 wire net223;
 wire net2230;
 wire net2231;
 wire net2232;
 wire net2233;
 wire net2234;
 wire net2235;
 wire net2236;
 wire net2237;
 wire net2238;
 wire net2239;
 wire net224;
 wire net2240;
 wire net2241;
 wire net2242;
 wire net2243;
 wire net2244;
 wire net2245;
 wire net2246;
 wire net2247;
 wire net2248;
 wire net2249;
 wire net225;
 wire net2250;
 wire net2251;
 wire net2252;
 wire net2253;
 wire net2254;
 wire net2255;
 wire net2256;
 wire net2257;
 wire net2258;
 wire net2259;
 wire net226;
 wire net2260;
 wire net2261;
 wire net2262;
 wire net2263;
 wire net2264;
 wire net2265;
 wire net2266;
 wire net2267;
 wire net2268;
 wire net2269;
 wire net227;
 wire net2270;
 wire net2271;
 wire net2272;
 wire net2273;
 wire net2274;
 wire net2275;
 wire net2276;
 wire net2277;
 wire net2278;
 wire net2279;
 wire net228;
 wire net2280;
 wire net2281;
 wire net2282;
 wire net2283;
 wire net2284;
 wire net2285;
 wire net2286;
 wire net2287;
 wire net2288;
 wire net2289;
 wire net229;
 wire net2290;
 wire net2291;
 wire net2292;
 wire net2293;
 wire net2294;
 wire net2295;
 wire net2296;
 wire net2297;
 wire net2298;
 wire net2299;
 wire net23;
 wire net230;
 wire net2300;
 wire net2301;
 wire net2302;
 wire net2303;
 wire net2304;
 wire net2305;
 wire net2306;
 wire net2307;
 wire net2308;
 wire net2309;
 wire net231;
 wire net2310;
 wire net2311;
 wire net2312;
 wire net2313;
 wire net2314;
 wire net2315;
 wire net2316;
 wire net2317;
 wire net2318;
 wire net2319;
 wire net232;
 wire net2320;
 wire net2321;
 wire net2322;
 wire net2323;
 wire net2324;
 wire net2325;
 wire net2326;
 wire net2327;
 wire net2328;
 wire net2329;
 wire net233;
 wire net2330;
 wire net2331;
 wire net2332;
 wire net2333;
 wire net2334;
 wire net2335;
 wire net2336;
 wire net2337;
 wire net2338;
 wire net2339;
 wire net234;
 wire net2340;
 wire net2341;
 wire net2342;
 wire net2343;
 wire net2344;
 wire net2345;
 wire net2346;
 wire net2347;
 wire net2348;
 wire net2349;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net24;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net25;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net26;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net27;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net28;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net29;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net3;
 wire net30;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net31;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net32;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net33;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net34;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net35;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net36;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net37;
 wire net370;
 wire net371;
 wire net372;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net38;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net39;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net4;
 wire net40;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net41;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net42;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net43;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net44;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net45;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net46;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net47;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net48;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net49;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net5;
 wire net50;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net51;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net52;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net53;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net54;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net55;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net56;
 wire net560;
 wire net561;
 wire net562;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net57;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net58;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net59;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net6;
 wire net60;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net61;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net62;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net63;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net64;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net65;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net66;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net67;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net68;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net69;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net7;
 wire net70;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net71;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net72;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net73;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net74;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net75;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net76;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net77;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net78;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net79;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net8;
 wire net80;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net81;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net82;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net83;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net84;
 wire net840;
 wire net841;
 wire net842;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net85;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net86;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net87;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net88;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net89;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net9;
 wire net90;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net91;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net92;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net93;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net94;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net95;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net96;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net97;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net98;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net99;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire \reg_blk_sel[0] ;
 wire \reg_blk_sel[1] ;
 wire \reg_blk_sel[2] ;
 wire \reg_blk_sel[3] ;
 wire \u_glbl_reg.cfg_gpio_dgmode ;
 wire \u_glbl_reg.cfg_mon_sel[0] ;
 wire \u_glbl_reg.cfg_mon_sel[1] ;
 wire \u_glbl_reg.cfg_mon_sel[2] ;
 wire \u_glbl_reg.cfg_mon_sel[3] ;
 wire \u_glbl_reg.cfg_multi_func_sel[0] ;
 wire \u_glbl_reg.cfg_multi_func_sel[10] ;
 wire \u_glbl_reg.cfg_multi_func_sel[11] ;
 wire \u_glbl_reg.cfg_multi_func_sel[12] ;
 wire \u_glbl_reg.cfg_multi_func_sel[13] ;
 wire \u_glbl_reg.cfg_multi_func_sel[14] ;
 wire \u_glbl_reg.cfg_multi_func_sel[15] ;
 wire \u_glbl_reg.cfg_multi_func_sel[16] ;
 wire \u_glbl_reg.cfg_multi_func_sel[17] ;
 wire \u_glbl_reg.cfg_multi_func_sel[18] ;
 wire \u_glbl_reg.cfg_multi_func_sel[19] ;
 wire \u_glbl_reg.cfg_multi_func_sel[1] ;
 wire \u_glbl_reg.cfg_multi_func_sel[20] ;
 wire \u_glbl_reg.cfg_multi_func_sel[21] ;
 wire \u_glbl_reg.cfg_multi_func_sel[22] ;
 wire \u_glbl_reg.cfg_multi_func_sel[23] ;
 wire \u_glbl_reg.cfg_multi_func_sel[24] ;
 wire \u_glbl_reg.cfg_multi_func_sel[25] ;
 wire \u_glbl_reg.cfg_multi_func_sel[26] ;
 wire \u_glbl_reg.cfg_multi_func_sel[27] ;
 wire \u_glbl_reg.cfg_multi_func_sel[28] ;
 wire \u_glbl_reg.cfg_multi_func_sel[29] ;
 wire \u_glbl_reg.cfg_multi_func_sel[2] ;
 wire \u_glbl_reg.cfg_multi_func_sel[30] ;
 wire \u_glbl_reg.cfg_multi_func_sel[31] ;
 wire \u_glbl_reg.cfg_multi_func_sel[3] ;
 wire \u_glbl_reg.cfg_multi_func_sel[4] ;
 wire \u_glbl_reg.cfg_multi_func_sel[5] ;
 wire \u_glbl_reg.cfg_multi_func_sel[6] ;
 wire \u_glbl_reg.cfg_multi_func_sel[7] ;
 wire \u_glbl_reg.cfg_multi_func_sel[8] ;
 wire \u_glbl_reg.cfg_multi_func_sel[9] ;
 wire \u_glbl_reg.cfg_ref_pll_div[0] ;
 wire \u_glbl_reg.cfg_ref_pll_div[1] ;
 wire \u_glbl_reg.cfg_ref_pll_div[2] ;
 wire \u_glbl_reg.cfg_rst_ctrl[0] ;
 wire \u_glbl_reg.cfg_rst_ctrl[10] ;
 wire \u_glbl_reg.cfg_rst_ctrl[11] ;
 wire \u_glbl_reg.cfg_rst_ctrl[12] ;
 wire \u_glbl_reg.cfg_rst_ctrl[13] ;
 wire \u_glbl_reg.cfg_rst_ctrl[14] ;
 wire \u_glbl_reg.cfg_rst_ctrl[15] ;
 wire \u_glbl_reg.cfg_rst_ctrl[16] ;
 wire \u_glbl_reg.cfg_rst_ctrl[17] ;
 wire \u_glbl_reg.cfg_rst_ctrl[18] ;
 wire \u_glbl_reg.cfg_rst_ctrl[19] ;
 wire \u_glbl_reg.cfg_rst_ctrl[1] ;
 wire \u_glbl_reg.cfg_rst_ctrl[20] ;
 wire \u_glbl_reg.cfg_rst_ctrl[21] ;
 wire \u_glbl_reg.cfg_rst_ctrl[22] ;
 wire \u_glbl_reg.cfg_rst_ctrl[23] ;
 wire \u_glbl_reg.cfg_rst_ctrl[24] ;
 wire \u_glbl_reg.cfg_rst_ctrl[25] ;
 wire \u_glbl_reg.cfg_rst_ctrl[26] ;
 wire \u_glbl_reg.cfg_rst_ctrl[27] ;
 wire \u_glbl_reg.cfg_rst_ctrl[28] ;
 wire \u_glbl_reg.cfg_rst_ctrl[29] ;
 wire \u_glbl_reg.cfg_rst_ctrl[2] ;
 wire \u_glbl_reg.cfg_rst_ctrl[30] ;
 wire \u_glbl_reg.cfg_rst_ctrl[31] ;
 wire \u_glbl_reg.cfg_rst_ctrl[3] ;
 wire \u_glbl_reg.cfg_rst_ctrl[4] ;
 wire \u_glbl_reg.cfg_rst_ctrl[5] ;
 wire \u_glbl_reg.cfg_rst_ctrl[6] ;
 wire \u_glbl_reg.cfg_rst_ctrl[7] ;
 wire \u_glbl_reg.cfg_rst_ctrl[8] ;
 wire \u_glbl_reg.cfg_rst_ctrl[9] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[0] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[1] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[2] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[3] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[4] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[5] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[6] ;
 wire \u_glbl_reg.cfg_rtc_clk_ctrl[7] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[0] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[1] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[2] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[3] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[4] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[5] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[6] ;
 wire \u_glbl_reg.cfg_usb_clk_ctrl[7] ;
 wire \u_glbl_reg.dbg_clk_div16 ;
 wire \u_glbl_reg.dbg_clk_mon ;
 wire \u_glbl_reg.dbg_clk_ref ;
 wire \u_glbl_reg.dbg_clk_ref_buf ;
 wire \u_glbl_reg.i2cm_intr_s ;
 wire \u_glbl_reg.i2cm_intr_ss ;
 wire \u_glbl_reg.ir_intr_s ;
 wire \u_glbl_reg.ir_intr_ss ;
 wire \u_glbl_reg.p_reset_n ;
 wire \u_glbl_reg.reg_12[0] ;
 wire \u_glbl_reg.reg_12[10] ;
 wire \u_glbl_reg.reg_12[11] ;
 wire \u_glbl_reg.reg_12[12] ;
 wire \u_glbl_reg.reg_12[13] ;
 wire \u_glbl_reg.reg_12[14] ;
 wire \u_glbl_reg.reg_12[15] ;
 wire \u_glbl_reg.reg_12[1] ;
 wire \u_glbl_reg.reg_12[2] ;
 wire \u_glbl_reg.reg_12[3] ;
 wire \u_glbl_reg.reg_12[4] ;
 wire \u_glbl_reg.reg_12[5] ;
 wire \u_glbl_reg.reg_12[6] ;
 wire \u_glbl_reg.reg_12[7] ;
 wire \u_glbl_reg.reg_12[8] ;
 wire \u_glbl_reg.reg_12[9] ;
 wire \u_glbl_reg.reg_15[0] ;
 wire \u_glbl_reg.reg_15[10] ;
 wire \u_glbl_reg.reg_15[11] ;
 wire \u_glbl_reg.reg_15[12] ;
 wire \u_glbl_reg.reg_15[13] ;
 wire \u_glbl_reg.reg_15[14] ;
 wire \u_glbl_reg.reg_15[15] ;
 wire \u_glbl_reg.reg_15[16] ;
 wire \u_glbl_reg.reg_15[17] ;
 wire \u_glbl_reg.reg_15[18] ;
 wire \u_glbl_reg.reg_15[19] ;
 wire \u_glbl_reg.reg_15[1] ;
 wire \u_glbl_reg.reg_15[20] ;
 wire \u_glbl_reg.reg_15[21] ;
 wire \u_glbl_reg.reg_15[22] ;
 wire \u_glbl_reg.reg_15[23] ;
 wire \u_glbl_reg.reg_15[24] ;
 wire \u_glbl_reg.reg_15[25] ;
 wire \u_glbl_reg.reg_15[26] ;
 wire \u_glbl_reg.reg_15[27] ;
 wire \u_glbl_reg.reg_15[28] ;
 wire \u_glbl_reg.reg_15[29] ;
 wire \u_glbl_reg.reg_15[2] ;
 wire \u_glbl_reg.reg_15[30] ;
 wire \u_glbl_reg.reg_15[31] ;
 wire \u_glbl_reg.reg_15[3] ;
 wire \u_glbl_reg.reg_15[4] ;
 wire \u_glbl_reg.reg_15[5] ;
 wire \u_glbl_reg.reg_15[6] ;
 wire \u_glbl_reg.reg_15[7] ;
 wire \u_glbl_reg.reg_15[8] ;
 wire \u_glbl_reg.reg_15[9] ;
 wire \u_glbl_reg.reg_16[0] ;
 wire \u_glbl_reg.reg_16[10] ;
 wire \u_glbl_reg.reg_16[11] ;
 wire \u_glbl_reg.reg_16[12] ;
 wire \u_glbl_reg.reg_16[13] ;
 wire \u_glbl_reg.reg_16[14] ;
 wire \u_glbl_reg.reg_16[15] ;
 wire \u_glbl_reg.reg_16[16] ;
 wire \u_glbl_reg.reg_16[17] ;
 wire \u_glbl_reg.reg_16[18] ;
 wire \u_glbl_reg.reg_16[19] ;
 wire \u_glbl_reg.reg_16[1] ;
 wire \u_glbl_reg.reg_16[20] ;
 wire \u_glbl_reg.reg_16[21] ;
 wire \u_glbl_reg.reg_16[22] ;
 wire \u_glbl_reg.reg_16[23] ;
 wire \u_glbl_reg.reg_16[24] ;
 wire \u_glbl_reg.reg_16[25] ;
 wire \u_glbl_reg.reg_16[26] ;
 wire \u_glbl_reg.reg_16[27] ;
 wire \u_glbl_reg.reg_16[28] ;
 wire \u_glbl_reg.reg_16[29] ;
 wire \u_glbl_reg.reg_16[2] ;
 wire \u_glbl_reg.reg_16[30] ;
 wire \u_glbl_reg.reg_16[31] ;
 wire \u_glbl_reg.reg_16[3] ;
 wire \u_glbl_reg.reg_16[4] ;
 wire \u_glbl_reg.reg_16[5] ;
 wire \u_glbl_reg.reg_16[6] ;
 wire \u_glbl_reg.reg_16[7] ;
 wire \u_glbl_reg.reg_16[8] ;
 wire \u_glbl_reg.reg_16[9] ;
 wire \u_glbl_reg.reg_17[0] ;
 wire \u_glbl_reg.reg_17[10] ;
 wire \u_glbl_reg.reg_17[11] ;
 wire \u_glbl_reg.reg_17[12] ;
 wire \u_glbl_reg.reg_17[13] ;
 wire \u_glbl_reg.reg_17[14] ;
 wire \u_glbl_reg.reg_17[15] ;
 wire \u_glbl_reg.reg_17[16] ;
 wire \u_glbl_reg.reg_17[17] ;
 wire \u_glbl_reg.reg_17[18] ;
 wire \u_glbl_reg.reg_17[19] ;
 wire \u_glbl_reg.reg_17[1] ;
 wire \u_glbl_reg.reg_17[20] ;
 wire \u_glbl_reg.reg_17[21] ;
 wire \u_glbl_reg.reg_17[22] ;
 wire \u_glbl_reg.reg_17[23] ;
 wire \u_glbl_reg.reg_17[24] ;
 wire \u_glbl_reg.reg_17[25] ;
 wire \u_glbl_reg.reg_17[26] ;
 wire \u_glbl_reg.reg_17[27] ;
 wire \u_glbl_reg.reg_17[28] ;
 wire \u_glbl_reg.reg_17[29] ;
 wire \u_glbl_reg.reg_17[2] ;
 wire \u_glbl_reg.reg_17[30] ;
 wire \u_glbl_reg.reg_17[31] ;
 wire \u_glbl_reg.reg_17[3] ;
 wire \u_glbl_reg.reg_17[4] ;
 wire \u_glbl_reg.reg_17[5] ;
 wire \u_glbl_reg.reg_17[6] ;
 wire \u_glbl_reg.reg_17[7] ;
 wire \u_glbl_reg.reg_17[8] ;
 wire \u_glbl_reg.reg_17[9] ;
 wire \u_glbl_reg.reg_18[0] ;
 wire \u_glbl_reg.reg_18[10] ;
 wire \u_glbl_reg.reg_18[11] ;
 wire \u_glbl_reg.reg_18[12] ;
 wire \u_glbl_reg.reg_18[13] ;
 wire \u_glbl_reg.reg_18[14] ;
 wire \u_glbl_reg.reg_18[15] ;
 wire \u_glbl_reg.reg_18[16] ;
 wire \u_glbl_reg.reg_18[17] ;
 wire \u_glbl_reg.reg_18[18] ;
 wire \u_glbl_reg.reg_18[19] ;
 wire \u_glbl_reg.reg_18[1] ;
 wire \u_glbl_reg.reg_18[20] ;
 wire \u_glbl_reg.reg_18[21] ;
 wire \u_glbl_reg.reg_18[22] ;
 wire \u_glbl_reg.reg_18[23] ;
 wire \u_glbl_reg.reg_18[24] ;
 wire \u_glbl_reg.reg_18[25] ;
 wire \u_glbl_reg.reg_18[26] ;
 wire \u_glbl_reg.reg_18[27] ;
 wire \u_glbl_reg.reg_18[28] ;
 wire \u_glbl_reg.reg_18[29] ;
 wire \u_glbl_reg.reg_18[2] ;
 wire \u_glbl_reg.reg_18[30] ;
 wire \u_glbl_reg.reg_18[31] ;
 wire \u_glbl_reg.reg_18[3] ;
 wire \u_glbl_reg.reg_18[4] ;
 wire \u_glbl_reg.reg_18[5] ;
 wire \u_glbl_reg.reg_18[6] ;
 wire \u_glbl_reg.reg_18[7] ;
 wire \u_glbl_reg.reg_18[8] ;
 wire \u_glbl_reg.reg_18[9] ;
 wire \u_glbl_reg.reg_19[0] ;
 wire \u_glbl_reg.reg_19[10] ;
 wire \u_glbl_reg.reg_19[11] ;
 wire \u_glbl_reg.reg_19[12] ;
 wire \u_glbl_reg.reg_19[13] ;
 wire \u_glbl_reg.reg_19[14] ;
 wire \u_glbl_reg.reg_19[15] ;
 wire \u_glbl_reg.reg_19[16] ;
 wire \u_glbl_reg.reg_19[17] ;
 wire \u_glbl_reg.reg_19[18] ;
 wire \u_glbl_reg.reg_19[19] ;
 wire \u_glbl_reg.reg_19[1] ;
 wire \u_glbl_reg.reg_19[20] ;
 wire \u_glbl_reg.reg_19[21] ;
 wire \u_glbl_reg.reg_19[22] ;
 wire \u_glbl_reg.reg_19[23] ;
 wire \u_glbl_reg.reg_19[24] ;
 wire \u_glbl_reg.reg_19[25] ;
 wire \u_glbl_reg.reg_19[26] ;
 wire \u_glbl_reg.reg_19[27] ;
 wire \u_glbl_reg.reg_19[28] ;
 wire \u_glbl_reg.reg_19[29] ;
 wire \u_glbl_reg.reg_19[2] ;
 wire \u_glbl_reg.reg_19[30] ;
 wire \u_glbl_reg.reg_19[31] ;
 wire \u_glbl_reg.reg_19[3] ;
 wire \u_glbl_reg.reg_19[4] ;
 wire \u_glbl_reg.reg_19[5] ;
 wire \u_glbl_reg.reg_19[6] ;
 wire \u_glbl_reg.reg_19[7] ;
 wire \u_glbl_reg.reg_19[8] ;
 wire \u_glbl_reg.reg_19[9] ;
 wire \u_glbl_reg.reg_20[0] ;
 wire \u_glbl_reg.reg_20[10] ;
 wire \u_glbl_reg.reg_20[11] ;
 wire \u_glbl_reg.reg_20[12] ;
 wire \u_glbl_reg.reg_20[13] ;
 wire \u_glbl_reg.reg_20[14] ;
 wire \u_glbl_reg.reg_20[15] ;
 wire \u_glbl_reg.reg_20[16] ;
 wire \u_glbl_reg.reg_20[17] ;
 wire \u_glbl_reg.reg_20[18] ;
 wire \u_glbl_reg.reg_20[19] ;
 wire \u_glbl_reg.reg_20[1] ;
 wire \u_glbl_reg.reg_20[20] ;
 wire \u_glbl_reg.reg_20[21] ;
 wire \u_glbl_reg.reg_20[22] ;
 wire \u_glbl_reg.reg_20[23] ;
 wire \u_glbl_reg.reg_20[24] ;
 wire \u_glbl_reg.reg_20[25] ;
 wire \u_glbl_reg.reg_20[26] ;
 wire \u_glbl_reg.reg_20[27] ;
 wire \u_glbl_reg.reg_20[28] ;
 wire \u_glbl_reg.reg_20[29] ;
 wire \u_glbl_reg.reg_20[2] ;
 wire \u_glbl_reg.reg_20[30] ;
 wire \u_glbl_reg.reg_20[31] ;
 wire \u_glbl_reg.reg_20[3] ;
 wire \u_glbl_reg.reg_20[4] ;
 wire \u_glbl_reg.reg_20[5] ;
 wire \u_glbl_reg.reg_20[6] ;
 wire \u_glbl_reg.reg_20[7] ;
 wire \u_glbl_reg.reg_20[8] ;
 wire \u_glbl_reg.reg_20[9] ;
 wire \u_glbl_reg.reg_21[0] ;
 wire \u_glbl_reg.reg_21[10] ;
 wire \u_glbl_reg.reg_21[11] ;
 wire \u_glbl_reg.reg_21[12] ;
 wire \u_glbl_reg.reg_21[13] ;
 wire \u_glbl_reg.reg_21[14] ;
 wire \u_glbl_reg.reg_21[15] ;
 wire \u_glbl_reg.reg_21[16] ;
 wire \u_glbl_reg.reg_21[17] ;
 wire \u_glbl_reg.reg_21[18] ;
 wire \u_glbl_reg.reg_21[19] ;
 wire \u_glbl_reg.reg_21[1] ;
 wire \u_glbl_reg.reg_21[20] ;
 wire \u_glbl_reg.reg_21[21] ;
 wire \u_glbl_reg.reg_21[22] ;
 wire \u_glbl_reg.reg_21[23] ;
 wire \u_glbl_reg.reg_21[24] ;
 wire \u_glbl_reg.reg_21[25] ;
 wire \u_glbl_reg.reg_21[26] ;
 wire \u_glbl_reg.reg_21[27] ;
 wire \u_glbl_reg.reg_21[28] ;
 wire \u_glbl_reg.reg_21[29] ;
 wire \u_glbl_reg.reg_21[2] ;
 wire \u_glbl_reg.reg_21[30] ;
 wire \u_glbl_reg.reg_21[31] ;
 wire \u_glbl_reg.reg_21[3] ;
 wire \u_glbl_reg.reg_21[4] ;
 wire \u_glbl_reg.reg_21[5] ;
 wire \u_glbl_reg.reg_21[6] ;
 wire \u_glbl_reg.reg_21[7] ;
 wire \u_glbl_reg.reg_21[8] ;
 wire \u_glbl_reg.reg_21[9] ;
 wire \u_glbl_reg.reg_22[0] ;
 wire \u_glbl_reg.reg_22[10] ;
 wire \u_glbl_reg.reg_22[11] ;
 wire \u_glbl_reg.reg_22[12] ;
 wire \u_glbl_reg.reg_22[13] ;
 wire \u_glbl_reg.reg_22[14] ;
 wire \u_glbl_reg.reg_22[15] ;
 wire \u_glbl_reg.reg_22[16] ;
 wire \u_glbl_reg.reg_22[17] ;
 wire \u_glbl_reg.reg_22[18] ;
 wire \u_glbl_reg.reg_22[19] ;
 wire \u_glbl_reg.reg_22[1] ;
 wire \u_glbl_reg.reg_22[20] ;
 wire \u_glbl_reg.reg_22[21] ;
 wire \u_glbl_reg.reg_22[22] ;
 wire \u_glbl_reg.reg_22[23] ;
 wire \u_glbl_reg.reg_22[24] ;
 wire \u_glbl_reg.reg_22[25] ;
 wire \u_glbl_reg.reg_22[26] ;
 wire \u_glbl_reg.reg_22[27] ;
 wire \u_glbl_reg.reg_22[28] ;
 wire \u_glbl_reg.reg_22[29] ;
 wire \u_glbl_reg.reg_22[2] ;
 wire \u_glbl_reg.reg_22[30] ;
 wire \u_glbl_reg.reg_22[31] ;
 wire \u_glbl_reg.reg_22[3] ;
 wire \u_glbl_reg.reg_22[4] ;
 wire \u_glbl_reg.reg_22[5] ;
 wire \u_glbl_reg.reg_22[6] ;
 wire \u_glbl_reg.reg_22[7] ;
 wire \u_glbl_reg.reg_22[8] ;
 wire \u_glbl_reg.reg_22[9] ;
 wire \u_glbl_reg.reg_23[0] ;
 wire \u_glbl_reg.reg_23[10] ;
 wire \u_glbl_reg.reg_23[11] ;
 wire \u_glbl_reg.reg_23[12] ;
 wire \u_glbl_reg.reg_23[13] ;
 wire \u_glbl_reg.reg_23[14] ;
 wire \u_glbl_reg.reg_23[15] ;
 wire \u_glbl_reg.reg_23[16] ;
 wire \u_glbl_reg.reg_23[17] ;
 wire \u_glbl_reg.reg_23[18] ;
 wire \u_glbl_reg.reg_23[19] ;
 wire \u_glbl_reg.reg_23[1] ;
 wire \u_glbl_reg.reg_23[20] ;
 wire \u_glbl_reg.reg_23[21] ;
 wire \u_glbl_reg.reg_23[22] ;
 wire \u_glbl_reg.reg_23[23] ;
 wire \u_glbl_reg.reg_23[24] ;
 wire \u_glbl_reg.reg_23[25] ;
 wire \u_glbl_reg.reg_23[26] ;
 wire \u_glbl_reg.reg_23[27] ;
 wire \u_glbl_reg.reg_23[28] ;
 wire \u_glbl_reg.reg_23[29] ;
 wire \u_glbl_reg.reg_23[2] ;
 wire \u_glbl_reg.reg_23[30] ;
 wire \u_glbl_reg.reg_23[31] ;
 wire \u_glbl_reg.reg_23[3] ;
 wire \u_glbl_reg.reg_23[4] ;
 wire \u_glbl_reg.reg_23[5] ;
 wire \u_glbl_reg.reg_23[6] ;
 wire \u_glbl_reg.reg_23[7] ;
 wire \u_glbl_reg.reg_23[8] ;
 wire \u_glbl_reg.reg_23[9] ;
 wire \u_glbl_reg.reg_2[0] ;
 wire \u_glbl_reg.reg_2[10] ;
 wire \u_glbl_reg.reg_2[11] ;
 wire \u_glbl_reg.reg_2[12] ;
 wire \u_glbl_reg.reg_2[13] ;
 wire \u_glbl_reg.reg_2[14] ;
 wire \u_glbl_reg.reg_2[15] ;
 wire \u_glbl_reg.reg_2[16] ;
 wire \u_glbl_reg.reg_2[17] ;
 wire \u_glbl_reg.reg_2[18] ;
 wire \u_glbl_reg.reg_2[19] ;
 wire \u_glbl_reg.reg_2[1] ;
 wire \u_glbl_reg.reg_2[20] ;
 wire \u_glbl_reg.reg_2[21] ;
 wire \u_glbl_reg.reg_2[22] ;
 wire \u_glbl_reg.reg_2[23] ;
 wire \u_glbl_reg.reg_2[24] ;
 wire \u_glbl_reg.reg_2[25] ;
 wire \u_glbl_reg.reg_2[26] ;
 wire \u_glbl_reg.reg_2[27] ;
 wire \u_glbl_reg.reg_2[28] ;
 wire \u_glbl_reg.reg_2[29] ;
 wire \u_glbl_reg.reg_2[2] ;
 wire \u_glbl_reg.reg_2[30] ;
 wire \u_glbl_reg.reg_2[31] ;
 wire \u_glbl_reg.reg_2[9] ;
 wire \u_glbl_reg.reg_3[0] ;
 wire \u_glbl_reg.reg_3[10] ;
 wire \u_glbl_reg.reg_3[11] ;
 wire \u_glbl_reg.reg_3[12] ;
 wire \u_glbl_reg.reg_3[13] ;
 wire \u_glbl_reg.reg_3[14] ;
 wire \u_glbl_reg.reg_3[15] ;
 wire \u_glbl_reg.reg_3[16] ;
 wire \u_glbl_reg.reg_3[17] ;
 wire \u_glbl_reg.reg_3[18] ;
 wire \u_glbl_reg.reg_3[19] ;
 wire \u_glbl_reg.reg_3[1] ;
 wire \u_glbl_reg.reg_3[20] ;
 wire \u_glbl_reg.reg_3[21] ;
 wire \u_glbl_reg.reg_3[22] ;
 wire \u_glbl_reg.reg_3[23] ;
 wire \u_glbl_reg.reg_3[24] ;
 wire \u_glbl_reg.reg_3[25] ;
 wire \u_glbl_reg.reg_3[26] ;
 wire \u_glbl_reg.reg_3[27] ;
 wire \u_glbl_reg.reg_3[28] ;
 wire \u_glbl_reg.reg_3[29] ;
 wire \u_glbl_reg.reg_3[2] ;
 wire \u_glbl_reg.reg_3[30] ;
 wire \u_glbl_reg.reg_3[31] ;
 wire \u_glbl_reg.reg_3[3] ;
 wire \u_glbl_reg.reg_3[4] ;
 wire \u_glbl_reg.reg_3[5] ;
 wire \u_glbl_reg.reg_3[6] ;
 wire \u_glbl_reg.reg_3[7] ;
 wire \u_glbl_reg.reg_3[8] ;
 wire \u_glbl_reg.reg_3[9] ;
 wire \u_glbl_reg.reg_6[16] ;
 wire \u_glbl_reg.reg_6[17] ;
 wire \u_glbl_reg.reg_6[18] ;
 wire \u_glbl_reg.reg_6[19] ;
 wire \u_glbl_reg.reg_6[20] ;
 wire \u_glbl_reg.reg_6[21] ;
 wire \u_glbl_reg.reg_6[22] ;
 wire \u_glbl_reg.reg_6[23] ;
 wire \u_glbl_reg.reg_6[24] ;
 wire \u_glbl_reg.reg_6[25] ;
 wire \u_glbl_reg.reg_6[26] ;
 wire \u_glbl_reg.reg_6[27] ;
 wire \u_glbl_reg.reg_6[28] ;
 wire \u_glbl_reg.reg_6[29] ;
 wire \u_glbl_reg.reg_6[30] ;
 wire \u_glbl_reg.reg_6[31] ;
 wire \u_glbl_reg.reg_7[10] ;
 wire \u_glbl_reg.reg_7[11] ;
 wire \u_glbl_reg.reg_7[12] ;
 wire \u_glbl_reg.reg_7[13] ;
 wire \u_glbl_reg.reg_7[14] ;
 wire \u_glbl_reg.reg_7[15] ;
 wire \u_glbl_reg.reg_7[16] ;
 wire \u_glbl_reg.reg_7[17] ;
 wire \u_glbl_reg.reg_7[18] ;
 wire \u_glbl_reg.reg_7[19] ;
 wire \u_glbl_reg.reg_7[20] ;
 wire \u_glbl_reg.reg_7[21] ;
 wire \u_glbl_reg.reg_7[22] ;
 wire \u_glbl_reg.reg_7[23] ;
 wire \u_glbl_reg.reg_7[24] ;
 wire \u_glbl_reg.reg_7[25] ;
 wire \u_glbl_reg.reg_7[26] ;
 wire \u_glbl_reg.reg_7[27] ;
 wire \u_glbl_reg.reg_7[28] ;
 wire \u_glbl_reg.reg_7[29] ;
 wire \u_glbl_reg.reg_7[30] ;
 wire \u_glbl_reg.reg_7[31] ;
 wire \u_glbl_reg.reg_7[4] ;
 wire \u_glbl_reg.reg_7[5] ;
 wire \u_glbl_reg.reg_7[6] ;
 wire \u_glbl_reg.reg_7[7] ;
 wire \u_glbl_reg.reg_7[8] ;
 wire \u_glbl_reg.reg_7[9] ;
 wire \u_glbl_reg.reg_ack ;
 wire \u_glbl_reg.reg_out[0] ;
 wire \u_glbl_reg.reg_out[10] ;
 wire \u_glbl_reg.reg_out[11] ;
 wire \u_glbl_reg.reg_out[12] ;
 wire \u_glbl_reg.reg_out[13] ;
 wire \u_glbl_reg.reg_out[14] ;
 wire \u_glbl_reg.reg_out[15] ;
 wire \u_glbl_reg.reg_out[16] ;
 wire \u_glbl_reg.reg_out[17] ;
 wire \u_glbl_reg.reg_out[18] ;
 wire \u_glbl_reg.reg_out[19] ;
 wire \u_glbl_reg.reg_out[1] ;
 wire \u_glbl_reg.reg_out[20] ;
 wire \u_glbl_reg.reg_out[21] ;
 wire \u_glbl_reg.reg_out[22] ;
 wire \u_glbl_reg.reg_out[23] ;
 wire \u_glbl_reg.reg_out[24] ;
 wire \u_glbl_reg.reg_out[25] ;
 wire \u_glbl_reg.reg_out[26] ;
 wire \u_glbl_reg.reg_out[27] ;
 wire \u_glbl_reg.reg_out[28] ;
 wire \u_glbl_reg.reg_out[29] ;
 wire \u_glbl_reg.reg_out[2] ;
 wire \u_glbl_reg.reg_out[30] ;
 wire \u_glbl_reg.reg_out[31] ;
 wire \u_glbl_reg.reg_out[3] ;
 wire \u_glbl_reg.reg_out[4] ;
 wire \u_glbl_reg.reg_out[5] ;
 wire \u_glbl_reg.reg_out[6] ;
 wire \u_glbl_reg.reg_out[7] ;
 wire \u_glbl_reg.reg_out[8] ;
 wire \u_glbl_reg.reg_out[9] ;
 wire \u_glbl_reg.reg_rdata[0] ;
 wire \u_glbl_reg.reg_rdata[10] ;
 wire \u_glbl_reg.reg_rdata[11] ;
 wire \u_glbl_reg.reg_rdata[12] ;
 wire \u_glbl_reg.reg_rdata[13] ;
 wire \u_glbl_reg.reg_rdata[14] ;
 wire \u_glbl_reg.reg_rdata[15] ;
 wire \u_glbl_reg.reg_rdata[16] ;
 wire \u_glbl_reg.reg_rdata[17] ;
 wire \u_glbl_reg.reg_rdata[18] ;
 wire \u_glbl_reg.reg_rdata[19] ;
 wire \u_glbl_reg.reg_rdata[1] ;
 wire \u_glbl_reg.reg_rdata[20] ;
 wire \u_glbl_reg.reg_rdata[21] ;
 wire \u_glbl_reg.reg_rdata[22] ;
 wire \u_glbl_reg.reg_rdata[23] ;
 wire \u_glbl_reg.reg_rdata[24] ;
 wire \u_glbl_reg.reg_rdata[25] ;
 wire \u_glbl_reg.reg_rdata[26] ;
 wire \u_glbl_reg.reg_rdata[27] ;
 wire \u_glbl_reg.reg_rdata[28] ;
 wire \u_glbl_reg.reg_rdata[29] ;
 wire \u_glbl_reg.reg_rdata[2] ;
 wire \u_glbl_reg.reg_rdata[30] ;
 wire \u_glbl_reg.reg_rdata[31] ;
 wire \u_glbl_reg.reg_rdata[3] ;
 wire \u_glbl_reg.reg_rdata[4] ;
 wire \u_glbl_reg.reg_rdata[5] ;
 wire \u_glbl_reg.reg_rdata[6] ;
 wire \u_glbl_reg.reg_rdata[7] ;
 wire \u_glbl_reg.reg_rdata[8] ;
 wire \u_glbl_reg.reg_rdata[9] ;
 wire \u_glbl_reg.rtc_clk_div ;
 wire \u_glbl_reg.rtc_clk_int ;
 wire \u_glbl_reg.rtc_intr_s ;
 wire \u_glbl_reg.rtc_intr_ss ;
 wire \u_glbl_reg.rtc_ref_clk ;
 wire \u_glbl_reg.rtc_ref_clk_int ;
 wire \u_glbl_reg.s_reset_n ;
 wire \u_glbl_reg.u_buf_cpu0_rst.X ;
 wire \u_glbl_reg.u_buf_cpu1_rst.X ;
 wire \u_glbl_reg.u_buf_cpu2_rst.X ;
 wire \u_glbl_reg.u_buf_cpu3_rst.X ;
 wire \u_glbl_reg.u_buf_uart0_rst.X ;
 wire \u_glbl_reg.u_buf_uart1_rst.X ;
 wire \u_glbl_reg.u_clkbuf_usb.A ;
 wire \u_glbl_reg.u_dbgclk.high_count[0] ;
 wire \u_glbl_reg.u_dbgclk.high_count[1] ;
 wire \u_glbl_reg.u_dbgclk.high_count[2] ;
 wire \u_glbl_reg.u_dbgclk.high_count[3] ;
 wire \u_glbl_reg.u_dbgclk.low_count[0] ;
 wire \u_glbl_reg.u_dbgclk.low_count[1] ;
 wire \u_glbl_reg.u_dbgclk.low_count[2] ;
 wire \u_glbl_reg.u_dbgclk.low_count[3] ;
 wire \u_glbl_reg.u_pll_ref_clk.high_count[0] ;
 wire \u_glbl_reg.u_pll_ref_clk.high_count[1] ;
 wire \u_glbl_reg.u_pll_ref_clk.high_count[2] ;
 wire \u_glbl_reg.u_pll_ref_clk.low_count[0] ;
 wire \u_glbl_reg.u_pll_ref_clk.low_count[1] ;
 wire \u_glbl_reg.u_pll_ref_clk.low_count[2] ;
 wire \u_glbl_reg.u_random.n0[0] ;
 wire \u_glbl_reg.u_random.n0[10] ;
 wire \u_glbl_reg.u_random.n0[11] ;
 wire \u_glbl_reg.u_random.n0[12] ;
 wire \u_glbl_reg.u_random.n0[13] ;
 wire \u_glbl_reg.u_random.n0[14] ;
 wire \u_glbl_reg.u_random.n0[15] ;
 wire \u_glbl_reg.u_random.n0[16] ;
 wire \u_glbl_reg.u_random.n0[17] ;
 wire \u_glbl_reg.u_random.n0[18] ;
 wire \u_glbl_reg.u_random.n0[19] ;
 wire \u_glbl_reg.u_random.n0[1] ;
 wire \u_glbl_reg.u_random.n0[20] ;
 wire \u_glbl_reg.u_random.n0[21] ;
 wire \u_glbl_reg.u_random.n0[22] ;
 wire \u_glbl_reg.u_random.n0[23] ;
 wire \u_glbl_reg.u_random.n0[24] ;
 wire \u_glbl_reg.u_random.n0[25] ;
 wire \u_glbl_reg.u_random.n0[26] ;
 wire \u_glbl_reg.u_random.n0[27] ;
 wire \u_glbl_reg.u_random.n0[28] ;
 wire \u_glbl_reg.u_random.n0[29] ;
 wire \u_glbl_reg.u_random.n0[2] ;
 wire \u_glbl_reg.u_random.n0[30] ;
 wire \u_glbl_reg.u_random.n0[31] ;
 wire \u_glbl_reg.u_random.n0[3] ;
 wire \u_glbl_reg.u_random.n0[4] ;
 wire \u_glbl_reg.u_random.n0[5] ;
 wire \u_glbl_reg.u_random.n0[6] ;
 wire \u_glbl_reg.u_random.n0[7] ;
 wire \u_glbl_reg.u_random.n0[8] ;
 wire \u_glbl_reg.u_random.n0[9] ;
 wire \u_glbl_reg.u_random.n1[0] ;
 wire \u_glbl_reg.u_random.n1[10] ;
 wire \u_glbl_reg.u_random.n1[11] ;
 wire \u_glbl_reg.u_random.n1[12] ;
 wire \u_glbl_reg.u_random.n1[13] ;
 wire \u_glbl_reg.u_random.n1[14] ;
 wire \u_glbl_reg.u_random.n1[15] ;
 wire \u_glbl_reg.u_random.n1[16] ;
 wire \u_glbl_reg.u_random.n1[17] ;
 wire \u_glbl_reg.u_random.n1[18] ;
 wire \u_glbl_reg.u_random.n1[19] ;
 wire \u_glbl_reg.u_random.n1[1] ;
 wire \u_glbl_reg.u_random.n1[20] ;
 wire \u_glbl_reg.u_random.n1[21] ;
 wire \u_glbl_reg.u_random.n1[22] ;
 wire \u_glbl_reg.u_random.n1[23] ;
 wire \u_glbl_reg.u_random.n1[24] ;
 wire \u_glbl_reg.u_random.n1[25] ;
 wire \u_glbl_reg.u_random.n1[26] ;
 wire \u_glbl_reg.u_random.n1[27] ;
 wire \u_glbl_reg.u_random.n1[28] ;
 wire \u_glbl_reg.u_random.n1[29] ;
 wire \u_glbl_reg.u_random.n1[2] ;
 wire \u_glbl_reg.u_random.n1[30] ;
 wire \u_glbl_reg.u_random.n1[31] ;
 wire \u_glbl_reg.u_random.n1[3] ;
 wire \u_glbl_reg.u_random.n1[4] ;
 wire \u_glbl_reg.u_random.n1[5] ;
 wire \u_glbl_reg.u_random.n1[6] ;
 wire \u_glbl_reg.u_random.n1[7] ;
 wire \u_glbl_reg.u_random.n1[8] ;
 wire \u_glbl_reg.u_random.n1[9] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[0] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[10] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[11] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[12] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[13] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[14] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[15] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[16] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[17] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[18] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[19] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[1] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[20] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[21] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[22] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[23] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[24] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[25] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[26] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[27] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[28] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[29] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[2] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[30] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[31] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[3] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[4] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[5] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[6] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[7] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[8] ;
 wire \u_glbl_reg.u_random.n1_plus_n0[9] ;
 wire \u_glbl_reg.u_random.s0[0] ;
 wire \u_glbl_reg.u_random.s0[10] ;
 wire \u_glbl_reg.u_random.s0[11] ;
 wire \u_glbl_reg.u_random.s0[12] ;
 wire \u_glbl_reg.u_random.s0[13] ;
 wire \u_glbl_reg.u_random.s0[14] ;
 wire \u_glbl_reg.u_random.s0[15] ;
 wire \u_glbl_reg.u_random.s0[16] ;
 wire \u_glbl_reg.u_random.s0[17] ;
 wire \u_glbl_reg.u_random.s0[18] ;
 wire \u_glbl_reg.u_random.s0[19] ;
 wire \u_glbl_reg.u_random.s0[1] ;
 wire \u_glbl_reg.u_random.s0[20] ;
 wire \u_glbl_reg.u_random.s0[21] ;
 wire \u_glbl_reg.u_random.s0[22] ;
 wire \u_glbl_reg.u_random.s0[23] ;
 wire \u_glbl_reg.u_random.s0[24] ;
 wire \u_glbl_reg.u_random.s0[25] ;
 wire \u_glbl_reg.u_random.s0[26] ;
 wire \u_glbl_reg.u_random.s0[27] ;
 wire \u_glbl_reg.u_random.s0[28] ;
 wire \u_glbl_reg.u_random.s0[29] ;
 wire \u_glbl_reg.u_random.s0[2] ;
 wire \u_glbl_reg.u_random.s0[30] ;
 wire \u_glbl_reg.u_random.s0[31] ;
 wire \u_glbl_reg.u_random.s0[3] ;
 wire \u_glbl_reg.u_random.s0[4] ;
 wire \u_glbl_reg.u_random.s0[5] ;
 wire \u_glbl_reg.u_random.s0[6] ;
 wire \u_glbl_reg.u_random.s0[7] ;
 wire \u_glbl_reg.u_random.s0[8] ;
 wire \u_glbl_reg.u_random.s0[9] ;
 wire \u_glbl_reg.u_random.s1[0] ;
 wire \u_glbl_reg.u_random.s1[10] ;
 wire \u_glbl_reg.u_random.s1[11] ;
 wire \u_glbl_reg.u_random.s1[12] ;
 wire \u_glbl_reg.u_random.s1[13] ;
 wire \u_glbl_reg.u_random.s1[14] ;
 wire \u_glbl_reg.u_random.s1[15] ;
 wire \u_glbl_reg.u_random.s1[16] ;
 wire \u_glbl_reg.u_random.s1[17] ;
 wire \u_glbl_reg.u_random.s1[18] ;
 wire \u_glbl_reg.u_random.s1[19] ;
 wire \u_glbl_reg.u_random.s1[1] ;
 wire \u_glbl_reg.u_random.s1[20] ;
 wire \u_glbl_reg.u_random.s1[21] ;
 wire \u_glbl_reg.u_random.s1[22] ;
 wire \u_glbl_reg.u_random.s1[23] ;
 wire \u_glbl_reg.u_random.s1[24] ;
 wire \u_glbl_reg.u_random.s1[25] ;
 wire \u_glbl_reg.u_random.s1[26] ;
 wire \u_glbl_reg.u_random.s1[27] ;
 wire \u_glbl_reg.u_random.s1[28] ;
 wire \u_glbl_reg.u_random.s1[29] ;
 wire \u_glbl_reg.u_random.s1[2] ;
 wire \u_glbl_reg.u_random.s1[30] ;
 wire \u_glbl_reg.u_random.s1[31] ;
 wire \u_glbl_reg.u_random.s1[3] ;
 wire \u_glbl_reg.u_random.s1[4] ;
 wire \u_glbl_reg.u_random.s1[5] ;
 wire \u_glbl_reg.u_random.s1[6] ;
 wire \u_glbl_reg.u_random.s1[7] ;
 wire \u_glbl_reg.u_random.s1[8] ;
 wire \u_glbl_reg.u_random.s1[9] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[0] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[10] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[11] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[12] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[13] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[14] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[15] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[16] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[17] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[18] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[19] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[1] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[20] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[21] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[22] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[23] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[24] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[25] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[26] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[27] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[28] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[29] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[2] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[30] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[31] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[3] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[4] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[5] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[6] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[7] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[8] ;
 wire \u_glbl_reg.u_random.s1_xor_s0[9] ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.data_out ;
 wire \u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.hware_req ;
 wire \u_glbl_reg.u_reg_1.flag ;
 wire \u_glbl_reg.u_rtcclk.high_count[0] ;
 wire \u_glbl_reg.u_rtcclk.high_count[1] ;
 wire \u_glbl_reg.u_rtcclk.high_count[2] ;
 wire \u_glbl_reg.u_rtcclk.high_count[3] ;
 wire \u_glbl_reg.u_rtcclk.high_count[4] ;
 wire \u_glbl_reg.u_rtcclk.low_count[0] ;
 wire \u_glbl_reg.u_rtcclk.low_count[1] ;
 wire \u_glbl_reg.u_rtcclk.low_count[2] ;
 wire \u_glbl_reg.u_rtcclk.low_count[3] ;
 wire \u_glbl_reg.u_rtcclk.low_count[4] ;
 wire \u_glbl_reg.u_usb_clk_sel.A0 ;
 wire \u_glbl_reg.u_usb_clk_sel.A1 ;
 wire \u_glbl_reg.u_usb_ref_clkbuf.A ;
 wire \u_glbl_reg.u_usbclk.high_count[0] ;
 wire \u_glbl_reg.u_usbclk.high_count[1] ;
 wire \u_glbl_reg.u_usbclk.high_count[2] ;
 wire \u_glbl_reg.u_usbclk.high_count[3] ;
 wire \u_glbl_reg.u_usbclk.high_count[4] ;
 wire \u_glbl_reg.u_usbclk.low_count[0] ;
 wire \u_glbl_reg.u_usbclk.low_count[1] ;
 wire \u_glbl_reg.u_usbclk.low_count[2] ;
 wire \u_glbl_reg.u_usbclk.low_count[3] ;
 wire \u_glbl_reg.u_usbclk.low_count[4] ;
 wire \u_glbl_reg.usb_intr_s ;
 wire \u_glbl_reg.usb_intr_ss ;
 wire \u_gpio.cfg_gpio_dir_sel[0] ;
 wire \u_gpio.cfg_gpio_dir_sel[10] ;
 wire \u_gpio.cfg_gpio_dir_sel[11] ;
 wire \u_gpio.cfg_gpio_dir_sel[12] ;
 wire \u_gpio.cfg_gpio_dir_sel[13] ;
 wire \u_gpio.cfg_gpio_dir_sel[14] ;
 wire \u_gpio.cfg_gpio_dir_sel[15] ;
 wire \u_gpio.cfg_gpio_dir_sel[16] ;
 wire \u_gpio.cfg_gpio_dir_sel[17] ;
 wire \u_gpio.cfg_gpio_dir_sel[18] ;
 wire \u_gpio.cfg_gpio_dir_sel[19] ;
 wire \u_gpio.cfg_gpio_dir_sel[1] ;
 wire \u_gpio.cfg_gpio_dir_sel[20] ;
 wire \u_gpio.cfg_gpio_dir_sel[21] ;
 wire \u_gpio.cfg_gpio_dir_sel[22] ;
 wire \u_gpio.cfg_gpio_dir_sel[23] ;
 wire \u_gpio.cfg_gpio_dir_sel[24] ;
 wire \u_gpio.cfg_gpio_dir_sel[25] ;
 wire \u_gpio.cfg_gpio_dir_sel[26] ;
 wire \u_gpio.cfg_gpio_dir_sel[27] ;
 wire \u_gpio.cfg_gpio_dir_sel[28] ;
 wire \u_gpio.cfg_gpio_dir_sel[29] ;
 wire \u_gpio.cfg_gpio_dir_sel[2] ;
 wire \u_gpio.cfg_gpio_dir_sel[30] ;
 wire \u_gpio.cfg_gpio_dir_sel[31] ;
 wire \u_gpio.cfg_gpio_dir_sel[3] ;
 wire \u_gpio.cfg_gpio_dir_sel[4] ;
 wire \u_gpio.cfg_gpio_dir_sel[5] ;
 wire \u_gpio.cfg_gpio_dir_sel[6] ;
 wire \u_gpio.cfg_gpio_dir_sel[7] ;
 wire \u_gpio.cfg_gpio_dir_sel[8] ;
 wire \u_gpio.cfg_gpio_dir_sel[9] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[0] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[10] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[11] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[12] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[13] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[14] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[15] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[16] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[17] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[18] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[19] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[1] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[20] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[21] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[22] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[23] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[24] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[25] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[26] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[27] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[28] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[29] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[2] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[30] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[31] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[3] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[4] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[5] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[6] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[7] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[8] ;
 wire \u_gpio.cfg_gpio_negedge_int_sel[9] ;
 wire \u_gpio.cfg_gpio_out_data[0] ;
 wire \u_gpio.cfg_gpio_out_data[10] ;
 wire \u_gpio.cfg_gpio_out_data[11] ;
 wire \u_gpio.cfg_gpio_out_data[12] ;
 wire \u_gpio.cfg_gpio_out_data[13] ;
 wire \u_gpio.cfg_gpio_out_data[14] ;
 wire \u_gpio.cfg_gpio_out_data[15] ;
 wire \u_gpio.cfg_gpio_out_data[16] ;
 wire \u_gpio.cfg_gpio_out_data[17] ;
 wire \u_gpio.cfg_gpio_out_data[18] ;
 wire \u_gpio.cfg_gpio_out_data[19] ;
 wire \u_gpio.cfg_gpio_out_data[1] ;
 wire \u_gpio.cfg_gpio_out_data[20] ;
 wire \u_gpio.cfg_gpio_out_data[21] ;
 wire \u_gpio.cfg_gpio_out_data[22] ;
 wire \u_gpio.cfg_gpio_out_data[23] ;
 wire \u_gpio.cfg_gpio_out_data[24] ;
 wire \u_gpio.cfg_gpio_out_data[25] ;
 wire \u_gpio.cfg_gpio_out_data[26] ;
 wire \u_gpio.cfg_gpio_out_data[27] ;
 wire \u_gpio.cfg_gpio_out_data[28] ;
 wire \u_gpio.cfg_gpio_out_data[29] ;
 wire \u_gpio.cfg_gpio_out_data[2] ;
 wire \u_gpio.cfg_gpio_out_data[30] ;
 wire \u_gpio.cfg_gpio_out_data[31] ;
 wire \u_gpio.cfg_gpio_out_data[3] ;
 wire \u_gpio.cfg_gpio_out_data[4] ;
 wire \u_gpio.cfg_gpio_out_data[5] ;
 wire \u_gpio.cfg_gpio_out_data[6] ;
 wire \u_gpio.cfg_gpio_out_data[7] ;
 wire \u_gpio.cfg_gpio_out_data[8] ;
 wire \u_gpio.cfg_gpio_out_data[9] ;
 wire \u_gpio.cfg_gpio_out_type[0] ;
 wire \u_gpio.cfg_gpio_out_type[10] ;
 wire \u_gpio.cfg_gpio_out_type[11] ;
 wire \u_gpio.cfg_gpio_out_type[12] ;
 wire \u_gpio.cfg_gpio_out_type[13] ;
 wire \u_gpio.cfg_gpio_out_type[14] ;
 wire \u_gpio.cfg_gpio_out_type[15] ;
 wire \u_gpio.cfg_gpio_out_type[16] ;
 wire \u_gpio.cfg_gpio_out_type[17] ;
 wire \u_gpio.cfg_gpio_out_type[18] ;
 wire \u_gpio.cfg_gpio_out_type[19] ;
 wire \u_gpio.cfg_gpio_out_type[1] ;
 wire \u_gpio.cfg_gpio_out_type[20] ;
 wire \u_gpio.cfg_gpio_out_type[21] ;
 wire \u_gpio.cfg_gpio_out_type[22] ;
 wire \u_gpio.cfg_gpio_out_type[23] ;
 wire \u_gpio.cfg_gpio_out_type[24] ;
 wire \u_gpio.cfg_gpio_out_type[25] ;
 wire \u_gpio.cfg_gpio_out_type[26] ;
 wire \u_gpio.cfg_gpio_out_type[27] ;
 wire \u_gpio.cfg_gpio_out_type[28] ;
 wire \u_gpio.cfg_gpio_out_type[29] ;
 wire \u_gpio.cfg_gpio_out_type[2] ;
 wire \u_gpio.cfg_gpio_out_type[30] ;
 wire \u_gpio.cfg_gpio_out_type[31] ;
 wire \u_gpio.cfg_gpio_out_type[3] ;
 wire \u_gpio.cfg_gpio_out_type[4] ;
 wire \u_gpio.cfg_gpio_out_type[5] ;
 wire \u_gpio.cfg_gpio_out_type[6] ;
 wire \u_gpio.cfg_gpio_out_type[7] ;
 wire \u_gpio.cfg_gpio_out_type[8] ;
 wire \u_gpio.cfg_gpio_out_type[9] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[0] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[10] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[11] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[12] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[13] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[14] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[15] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[16] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[17] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[18] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[19] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[1] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[20] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[21] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[22] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[23] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[24] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[25] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[26] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[27] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[28] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[29] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[2] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[30] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[31] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[3] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[4] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[5] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[6] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[7] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[8] ;
 wire \u_gpio.cfg_gpio_posedge_int_sel[9] ;
 wire \u_gpio.pulse_1us ;
 wire \u_gpio.reg_ack ;
 wire \u_gpio.reg_rdata[0] ;
 wire \u_gpio.reg_rdata[10] ;
 wire \u_gpio.reg_rdata[11] ;
 wire \u_gpio.reg_rdata[12] ;
 wire \u_gpio.reg_rdata[13] ;
 wire \u_gpio.reg_rdata[14] ;
 wire \u_gpio.reg_rdata[15] ;
 wire \u_gpio.reg_rdata[16] ;
 wire \u_gpio.reg_rdata[17] ;
 wire \u_gpio.reg_rdata[18] ;
 wire \u_gpio.reg_rdata[19] ;
 wire \u_gpio.reg_rdata[1] ;
 wire \u_gpio.reg_rdata[20] ;
 wire \u_gpio.reg_rdata[21] ;
 wire \u_gpio.reg_rdata[22] ;
 wire \u_gpio.reg_rdata[23] ;
 wire \u_gpio.reg_rdata[24] ;
 wire \u_gpio.reg_rdata[25] ;
 wire \u_gpio.reg_rdata[26] ;
 wire \u_gpio.reg_rdata[27] ;
 wire \u_gpio.reg_rdata[28] ;
 wire \u_gpio.reg_rdata[29] ;
 wire \u_gpio.reg_rdata[2] ;
 wire \u_gpio.reg_rdata[30] ;
 wire \u_gpio.reg_rdata[31] ;
 wire \u_gpio.reg_rdata[3] ;
 wire \u_gpio.reg_rdata[4] ;
 wire \u_gpio.reg_rdata[5] ;
 wire \u_gpio.reg_rdata[6] ;
 wire \u_gpio.reg_rdata[7] ;
 wire \u_gpio.reg_rdata[8] ;
 wire \u_gpio.reg_rdata[9] ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[0].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[10].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[11].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[12].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[13].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[14].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[15].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[16].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[17].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[18].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[19].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[1].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[20].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[21].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[22].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[24].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[25].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[26].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[27].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[28].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[29].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[2].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[30].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[31].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[3].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[4].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[8].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_out ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_reg ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_ss[0] ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_ss[1] ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_ss[2] ;
 wire \u_gpio.u_bit[9].u_dglitch.gpio_ss[3] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[0] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[10] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[11] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[12] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[13] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[14] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[15] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[16] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[17] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[18] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[19] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[1] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[20] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[21] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[22] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[23] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[24] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[25] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[26] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[27] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[28] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[29] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[2] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[30] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[31] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[3] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[4] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[5] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[6] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[7] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[8] ;
 wire \u_gpio.u_reg.cfg_gpio_int_mask[9] ;
 wire \u_gpio.u_reg.reg_out[0] ;
 wire \u_gpio.u_reg.reg_out[10] ;
 wire \u_gpio.u_reg.reg_out[11] ;
 wire \u_gpio.u_reg.reg_out[12] ;
 wire \u_gpio.u_reg.reg_out[13] ;
 wire \u_gpio.u_reg.reg_out[14] ;
 wire \u_gpio.u_reg.reg_out[15] ;
 wire \u_gpio.u_reg.reg_out[16] ;
 wire \u_gpio.u_reg.reg_out[17] ;
 wire \u_gpio.u_reg.reg_out[18] ;
 wire \u_gpio.u_reg.reg_out[19] ;
 wire \u_gpio.u_reg.reg_out[1] ;
 wire \u_gpio.u_reg.reg_out[20] ;
 wire \u_gpio.u_reg.reg_out[21] ;
 wire \u_gpio.u_reg.reg_out[22] ;
 wire \u_gpio.u_reg.reg_out[23] ;
 wire \u_gpio.u_reg.reg_out[24] ;
 wire \u_gpio.u_reg.reg_out[25] ;
 wire \u_gpio.u_reg.reg_out[26] ;
 wire \u_gpio.u_reg.reg_out[27] ;
 wire \u_gpio.u_reg.reg_out[28] ;
 wire \u_gpio.u_reg.reg_out[29] ;
 wire \u_gpio.u_reg.reg_out[2] ;
 wire \u_gpio.u_reg.reg_out[30] ;
 wire \u_gpio.u_reg.reg_out[31] ;
 wire \u_gpio.u_reg.reg_out[3] ;
 wire \u_gpio.u_reg.reg_out[4] ;
 wire \u_gpio.u_reg.reg_out[5] ;
 wire \u_gpio.u_reg.reg_out[6] ;
 wire \u_gpio.u_reg.reg_out[7] ;
 wire \u_gpio.u_reg.reg_out[8] ;
 wire \u_gpio.u_reg.reg_out[9] ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.hware_req ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.data_out ;
 wire \u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.hware_req ;
 wire \u_prst_sync.in_data_2s ;
 wire \u_prst_sync.in_data_s ;
 wire \u_pwm.blk_sel[0] ;
 wire \u_pwm.blk_sel[1] ;
 wire \u_pwm.blk_sel[2] ;
 wire \u_pwm.reg_ack_glbl ;
 wire \u_pwm.reg_ack_pwm0 ;
 wire \u_pwm.reg_ack_pwm1 ;
 wire \u_pwm.reg_ack_pwm2 ;
 wire \u_pwm.reg_rdata_glbl[0] ;
 wire \u_pwm.reg_rdata_glbl[10] ;
 wire \u_pwm.reg_rdata_glbl[16] ;
 wire \u_pwm.reg_rdata_glbl[17] ;
 wire \u_pwm.reg_rdata_glbl[18] ;
 wire \u_pwm.reg_rdata_glbl[1] ;
 wire \u_pwm.reg_rdata_glbl[2] ;
 wire \u_pwm.reg_rdata_glbl[3] ;
 wire \u_pwm.reg_rdata_glbl[4] ;
 wire \u_pwm.reg_rdata_glbl[5] ;
 wire \u_pwm.reg_rdata_glbl[8] ;
 wire \u_pwm.reg_rdata_glbl[9] ;
 wire \u_pwm.reg_rdata_pwm0[0] ;
 wire \u_pwm.reg_rdata_pwm0[10] ;
 wire \u_pwm.reg_rdata_pwm0[11] ;
 wire \u_pwm.reg_rdata_pwm0[12] ;
 wire \u_pwm.reg_rdata_pwm0[13] ;
 wire \u_pwm.reg_rdata_pwm0[14] ;
 wire \u_pwm.reg_rdata_pwm0[15] ;
 wire \u_pwm.reg_rdata_pwm0[16] ;
 wire \u_pwm.reg_rdata_pwm0[17] ;
 wire \u_pwm.reg_rdata_pwm0[18] ;
 wire \u_pwm.reg_rdata_pwm0[19] ;
 wire \u_pwm.reg_rdata_pwm0[1] ;
 wire \u_pwm.reg_rdata_pwm0[20] ;
 wire \u_pwm.reg_rdata_pwm0[21] ;
 wire \u_pwm.reg_rdata_pwm0[22] ;
 wire \u_pwm.reg_rdata_pwm0[23] ;
 wire \u_pwm.reg_rdata_pwm0[24] ;
 wire \u_pwm.reg_rdata_pwm0[25] ;
 wire \u_pwm.reg_rdata_pwm0[26] ;
 wire \u_pwm.reg_rdata_pwm0[27] ;
 wire \u_pwm.reg_rdata_pwm0[28] ;
 wire \u_pwm.reg_rdata_pwm0[29] ;
 wire \u_pwm.reg_rdata_pwm0[2] ;
 wire \u_pwm.reg_rdata_pwm0[30] ;
 wire \u_pwm.reg_rdata_pwm0[31] ;
 wire \u_pwm.reg_rdata_pwm0[3] ;
 wire \u_pwm.reg_rdata_pwm0[4] ;
 wire \u_pwm.reg_rdata_pwm0[5] ;
 wire \u_pwm.reg_rdata_pwm0[6] ;
 wire \u_pwm.reg_rdata_pwm0[7] ;
 wire \u_pwm.reg_rdata_pwm0[8] ;
 wire \u_pwm.reg_rdata_pwm0[9] ;
 wire \u_pwm.reg_rdata_pwm1[0] ;
 wire \u_pwm.reg_rdata_pwm1[10] ;
 wire \u_pwm.reg_rdata_pwm1[11] ;
 wire \u_pwm.reg_rdata_pwm1[12] ;
 wire \u_pwm.reg_rdata_pwm1[13] ;
 wire \u_pwm.reg_rdata_pwm1[14] ;
 wire \u_pwm.reg_rdata_pwm1[15] ;
 wire \u_pwm.reg_rdata_pwm1[16] ;
 wire \u_pwm.reg_rdata_pwm1[17] ;
 wire \u_pwm.reg_rdata_pwm1[18] ;
 wire \u_pwm.reg_rdata_pwm1[19] ;
 wire \u_pwm.reg_rdata_pwm1[1] ;
 wire \u_pwm.reg_rdata_pwm1[20] ;
 wire \u_pwm.reg_rdata_pwm1[21] ;
 wire \u_pwm.reg_rdata_pwm1[22] ;
 wire \u_pwm.reg_rdata_pwm1[23] ;
 wire \u_pwm.reg_rdata_pwm1[24] ;
 wire \u_pwm.reg_rdata_pwm1[25] ;
 wire \u_pwm.reg_rdata_pwm1[26] ;
 wire \u_pwm.reg_rdata_pwm1[27] ;
 wire \u_pwm.reg_rdata_pwm1[28] ;
 wire \u_pwm.reg_rdata_pwm1[29] ;
 wire \u_pwm.reg_rdata_pwm1[2] ;
 wire \u_pwm.reg_rdata_pwm1[30] ;
 wire \u_pwm.reg_rdata_pwm1[31] ;
 wire \u_pwm.reg_rdata_pwm1[3] ;
 wire \u_pwm.reg_rdata_pwm1[4] ;
 wire \u_pwm.reg_rdata_pwm1[5] ;
 wire \u_pwm.reg_rdata_pwm1[6] ;
 wire \u_pwm.reg_rdata_pwm1[7] ;
 wire \u_pwm.reg_rdata_pwm1[8] ;
 wire \u_pwm.reg_rdata_pwm1[9] ;
 wire \u_pwm.reg_rdata_pwm2[0] ;
 wire \u_pwm.reg_rdata_pwm2[10] ;
 wire \u_pwm.reg_rdata_pwm2[11] ;
 wire \u_pwm.reg_rdata_pwm2[12] ;
 wire \u_pwm.reg_rdata_pwm2[13] ;
 wire \u_pwm.reg_rdata_pwm2[14] ;
 wire \u_pwm.reg_rdata_pwm2[15] ;
 wire \u_pwm.reg_rdata_pwm2[16] ;
 wire \u_pwm.reg_rdata_pwm2[17] ;
 wire \u_pwm.reg_rdata_pwm2[18] ;
 wire \u_pwm.reg_rdata_pwm2[19] ;
 wire \u_pwm.reg_rdata_pwm2[1] ;
 wire \u_pwm.reg_rdata_pwm2[20] ;
 wire \u_pwm.reg_rdata_pwm2[21] ;
 wire \u_pwm.reg_rdata_pwm2[22] ;
 wire \u_pwm.reg_rdata_pwm2[23] ;
 wire \u_pwm.reg_rdata_pwm2[24] ;
 wire \u_pwm.reg_rdata_pwm2[25] ;
 wire \u_pwm.reg_rdata_pwm2[26] ;
 wire \u_pwm.reg_rdata_pwm2[27] ;
 wire \u_pwm.reg_rdata_pwm2[28] ;
 wire \u_pwm.reg_rdata_pwm2[29] ;
 wire \u_pwm.reg_rdata_pwm2[2] ;
 wire \u_pwm.reg_rdata_pwm2[30] ;
 wire \u_pwm.reg_rdata_pwm2[31] ;
 wire \u_pwm.reg_rdata_pwm2[3] ;
 wire \u_pwm.reg_rdata_pwm2[4] ;
 wire \u_pwm.reg_rdata_pwm2[5] ;
 wire \u_pwm.reg_rdata_pwm2[6] ;
 wire \u_pwm.reg_rdata_pwm2[7] ;
 wire \u_pwm.reg_rdata_pwm2[8] ;
 wire \u_pwm.reg_rdata_pwm2[9] ;
 wire \u_pwm.u_glbl_reg.reg_out[0] ;
 wire \u_pwm.u_glbl_reg.reg_out[10] ;
 wire \u_pwm.u_glbl_reg.reg_out[16] ;
 wire \u_pwm.u_glbl_reg.reg_out[17] ;
 wire \u_pwm.u_glbl_reg.reg_out[18] ;
 wire \u_pwm.u_glbl_reg.reg_out[1] ;
 wire \u_pwm.u_glbl_reg.reg_out[2] ;
 wire \u_pwm.u_glbl_reg.reg_out[3] ;
 wire \u_pwm.u_glbl_reg.reg_out[4] ;
 wire \u_pwm.u_glbl_reg.reg_out[5] ;
 wire \u_pwm.u_glbl_reg.reg_out[8] ;
 wire \u_pwm.u_glbl_reg.reg_out[9] ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[1].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[3].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[4].u_bit_reg.data_out ;
 wire \u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[5].u_bit_reg.data_out ;
 wire \u_pwm.u_pwm_0.cfg_comp0_center ;
 wire \u_pwm.u_pwm_0.cfg_comp1_center ;
 wire \u_pwm.u_pwm_0.cfg_comp2_center ;
 wire \u_pwm.u_pwm_0.cfg_comp3_center ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[10] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[11] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[12] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[13] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[14] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[15] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[4] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[5] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[6] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[7] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[8] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp0[9] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[10] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[11] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[12] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[13] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[14] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[15] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[4] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[5] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[6] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[7] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[8] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp1[9] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[10] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[11] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[12] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[13] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[14] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[15] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[4] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[5] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[6] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[7] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[8] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp2[9] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[10] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[11] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[12] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[13] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[14] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[15] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[4] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[5] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[6] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[7] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[8] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_comp3[9] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_dupdate ;
 wire \u_pwm.u_pwm_0.cfg_pwm_enb ;
 wire \u_pwm.u_pwm_0.cfg_pwm_gpio_edge ;
 wire \u_pwm.u_pwm_0.cfg_pwm_gpio_enb ;
 wire \u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_gpio_sel[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_gpio_sel[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_hold ;
 wire \u_pwm.u_pwm_0.cfg_pwm_inv ;
 wire \u_pwm.u_pwm_0.cfg_pwm_mode[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_mode[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_oneshot ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[10] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[11] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[12] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[13] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[14] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[15] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[4] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[5] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[6] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[7] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[8] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_period[9] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_run ;
 wire \u_pwm.u_pwm_0.cfg_pwm_scale[0] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_scale[1] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_scale[2] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_scale[3] ;
 wire \u_pwm.u_pwm_0.cfg_pwm_zeropd ;
 wire \u_pwm.u_pwm_0.gpio_tgr ;
 wire \u_pwm.u_pwm_0.u_pwm.gpio_l ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[15] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_ovflow ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_ovflow_l ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[11] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[13] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[14] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[3] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[5] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[7] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_scnt[9] ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_wfm_i ;
 wire \u_pwm.u_pwm_0.u_pwm.pwm_wfm_r ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[0] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[10] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[11] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[12] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[13] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[14] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[15] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[16] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[17] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[18] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[19] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[1] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[20] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[21] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[22] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[23] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[24] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[25] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[26] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[27] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[28] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[29] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[2] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[30] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[31] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[3] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[4] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[5] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[6] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[7] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[8] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_0[9] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[0] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[10] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[11] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[12] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[13] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[14] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[15] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[16] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[17] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[18] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[19] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[1] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[20] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[21] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[22] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[23] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[24] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[25] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[26] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[27] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[28] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[29] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[2] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[30] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[31] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[3] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[4] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[5] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[6] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[7] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[8] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_1[9] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[0] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[10] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[11] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[12] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[13] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[14] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[15] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[16] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[17] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[18] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[19] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[1] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[20] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[21] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[22] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[23] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[24] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[25] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[26] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[27] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[28] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[29] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[2] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[30] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[31] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[3] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[4] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[5] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[6] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[7] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[8] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_2[9] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[0] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[10] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[11] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[12] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[13] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[14] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[15] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[16] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[17] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[18] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[19] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[1] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[20] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[21] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[22] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[23] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[24] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[25] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[26] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[27] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[28] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[29] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[2] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[30] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[31] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[3] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[4] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[5] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[6] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[7] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[8] ;
 wire \u_pwm.u_pwm_0.u_reg.reg_out[9] ;
 wire \u_pwm.u_pwm_1.cfg_comp0_center ;
 wire \u_pwm.u_pwm_1.cfg_comp1_center ;
 wire \u_pwm.u_pwm_1.cfg_comp2_center ;
 wire \u_pwm.u_pwm_1.cfg_comp3_center ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[10] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[11] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[12] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[13] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[14] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[15] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[4] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[5] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[6] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[7] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[8] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp0[9] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[10] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[11] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[12] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[13] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[14] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[15] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[4] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[5] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[6] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[7] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[8] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp1[9] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[10] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[11] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[12] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[13] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[14] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[15] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[4] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[5] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[6] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[7] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[8] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp2[9] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[10] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[11] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[12] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[13] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[14] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[15] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[4] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[5] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[6] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[7] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[8] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_comp3[9] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_dupdate ;
 wire \u_pwm.u_pwm_1.cfg_pwm_enb ;
 wire \u_pwm.u_pwm_1.cfg_pwm_gpio_edge ;
 wire \u_pwm.u_pwm_1.cfg_pwm_gpio_enb ;
 wire \u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_gpio_sel[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_gpio_sel[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_hold ;
 wire \u_pwm.u_pwm_1.cfg_pwm_inv ;
 wire \u_pwm.u_pwm_1.cfg_pwm_mode[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_mode[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_oneshot ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[10] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[11] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[12] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[13] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[14] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[15] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[4] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[5] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[6] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[7] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[8] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_period[9] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_run ;
 wire \u_pwm.u_pwm_1.cfg_pwm_scale[0] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_scale[1] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_scale[2] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_scale[3] ;
 wire \u_pwm.u_pwm_1.cfg_pwm_zeropd ;
 wire \u_pwm.u_pwm_1.gpio_tgr ;
 wire \u_pwm.u_pwm_1.u_pwm.gpio_l ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[5] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_ovflow ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_ovflow_l ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[11] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[13] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[14] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[3] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[5] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[7] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_scnt[9] ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_wfm_i ;
 wire \u_pwm.u_pwm_1.u_pwm.pwm_wfm_r ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[0] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[10] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[11] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[12] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[13] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[14] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[15] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[16] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[17] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[18] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[19] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[1] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[20] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[21] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[22] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[23] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[24] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[25] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[26] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[27] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[28] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[29] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[2] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[30] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[31] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[3] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[4] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[5] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[6] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[7] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[8] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_0[9] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[0] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[10] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[11] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[12] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[13] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[14] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[15] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[16] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[17] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[18] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[19] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[1] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[20] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[21] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[22] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[23] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[24] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[25] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[26] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[27] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[28] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[29] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[2] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[30] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[31] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[3] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[4] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[5] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[6] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[7] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[8] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_1[9] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[0] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[10] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[11] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[12] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[13] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[14] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[15] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[16] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[17] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[18] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[19] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[1] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[20] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[21] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[22] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[23] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[24] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[25] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[26] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[27] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[28] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[29] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[2] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[30] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[31] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[3] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[4] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[5] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[6] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[7] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[8] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_2[9] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[0] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[10] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[11] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[12] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[13] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[14] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[15] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[16] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[17] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[18] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[19] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[1] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[20] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[21] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[22] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[23] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[24] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[25] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[26] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[27] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[28] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[29] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[2] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[30] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[31] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[3] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[4] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[5] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[6] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[7] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[8] ;
 wire \u_pwm.u_pwm_1.u_reg.reg_out[9] ;
 wire \u_pwm.u_pwm_2.cfg_comp0_center ;
 wire \u_pwm.u_pwm_2.cfg_comp1_center ;
 wire \u_pwm.u_pwm_2.cfg_comp2_center ;
 wire \u_pwm.u_pwm_2.cfg_comp3_center ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[10] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[11] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[12] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[13] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[14] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[15] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[4] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[5] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[6] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[7] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[8] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp0[9] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[10] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[11] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[12] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[13] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[14] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[15] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[4] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[5] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[6] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[7] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[8] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp1[9] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[10] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[11] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[12] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[13] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[14] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[15] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[4] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[5] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[6] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[7] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[8] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp2[9] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[10] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[11] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[12] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[13] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[14] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[15] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[4] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[5] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[6] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[7] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[8] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_comp3[9] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_dupdate ;
 wire \u_pwm.u_pwm_2.cfg_pwm_enb ;
 wire \u_pwm.u_pwm_2.cfg_pwm_gpio_edge ;
 wire \u_pwm.u_pwm_2.cfg_pwm_gpio_enb ;
 wire \u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_gpio_sel[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_hold ;
 wire \u_pwm.u_pwm_2.cfg_pwm_inv ;
 wire \u_pwm.u_pwm_2.cfg_pwm_mode[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_mode[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_oneshot ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[10] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[11] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[12] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[13] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[14] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[15] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[4] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[5] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[6] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[7] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[8] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_period[9] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_run ;
 wire \u_pwm.u_pwm_2.cfg_pwm_scale[0] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_scale[1] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_scale[2] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_scale[3] ;
 wire \u_pwm.u_pwm_2.cfg_pwm_zeropd ;
 wire \u_pwm.u_pwm_2.gpio_tgr ;
 wire \u_pwm.u_pwm_2.u_pwm.gpio_l ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[10] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[14] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[15] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_ovflow ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_ovflow_l ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[11] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[13] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[14] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[3] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[5] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[7] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_scnt[9] ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_wfm_i ;
 wire \u_pwm.u_pwm_2.u_pwm.pwm_wfm_r ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[0] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[10] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[11] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[12] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[13] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[14] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[15] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[16] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[17] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[18] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[19] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[1] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[20] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[21] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[22] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[23] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[24] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[25] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[26] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[27] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[28] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[29] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[2] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[30] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[31] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[3] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[4] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[5] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[6] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[7] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[8] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_0[9] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[0] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[10] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[11] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[12] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[13] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[14] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[15] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[16] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[17] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[18] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[19] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[1] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[20] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[21] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[22] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[23] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[24] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[25] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[26] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[27] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[28] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[29] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[2] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[30] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[31] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[3] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[4] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[5] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[6] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[7] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[8] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_1[9] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[0] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[10] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[11] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[12] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[13] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[14] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[15] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[16] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[17] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[18] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[19] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[1] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[20] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[21] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[22] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[23] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[24] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[25] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[26] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[27] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[28] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[29] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[2] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[30] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[31] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[3] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[4] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[5] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[6] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[7] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[8] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_2[9] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[0] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[10] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[11] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[12] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[13] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[14] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[15] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[16] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[17] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[18] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[19] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[1] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[20] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[21] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[22] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[23] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[24] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[25] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[26] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[27] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[28] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[29] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[2] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[30] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[31] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[3] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[4] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[5] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[6] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[7] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[8] ;
 wire \u_pwm.u_pwm_2.u_reg.reg_out[9] ;
 wire \u_rst_sync.in_data_2s ;
 wire \u_rst_sync.in_data_s ;
 wire \u_semaphore.reg_0[0] ;
 wire \u_semaphore.reg_0[10] ;
 wire \u_semaphore.reg_0[11] ;
 wire \u_semaphore.reg_0[12] ;
 wire \u_semaphore.reg_0[13] ;
 wire \u_semaphore.reg_0[14] ;
 wire \u_semaphore.reg_0[15] ;
 wire \u_semaphore.reg_0[1] ;
 wire \u_semaphore.reg_0[2] ;
 wire \u_semaphore.reg_0[3] ;
 wire \u_semaphore.reg_0[4] ;
 wire \u_semaphore.reg_0[5] ;
 wire \u_semaphore.reg_0[6] ;
 wire \u_semaphore.reg_0[7] ;
 wire \u_semaphore.reg_0[8] ;
 wire \u_semaphore.reg_0[9] ;
 wire \u_semaphore.reg_ack ;
 wire \u_semaphore.reg_out[0] ;
 wire \u_semaphore.reg_out[10] ;
 wire \u_semaphore.reg_out[11] ;
 wire \u_semaphore.reg_out[12] ;
 wire \u_semaphore.reg_out[13] ;
 wire \u_semaphore.reg_out[14] ;
 wire \u_semaphore.reg_out[15] ;
 wire \u_semaphore.reg_out[1] ;
 wire \u_semaphore.reg_out[2] ;
 wire \u_semaphore.reg_out[3] ;
 wire \u_semaphore.reg_out[4] ;
 wire \u_semaphore.reg_out[5] ;
 wire \u_semaphore.reg_out[6] ;
 wire \u_semaphore.reg_out[7] ;
 wire \u_semaphore.reg_out[8] ;
 wire \u_semaphore.reg_out[9] ;
 wire \u_semaphore.reg_rdata[0] ;
 wire \u_semaphore.reg_rdata[10] ;
 wire \u_semaphore.reg_rdata[11] ;
 wire \u_semaphore.reg_rdata[12] ;
 wire \u_semaphore.reg_rdata[13] ;
 wire \u_semaphore.reg_rdata[14] ;
 wire \u_semaphore.reg_rdata[15] ;
 wire \u_semaphore.reg_rdata[1] ;
 wire \u_semaphore.reg_rdata[2] ;
 wire \u_semaphore.reg_rdata[3] ;
 wire \u_semaphore.reg_rdata[4] ;
 wire \u_semaphore.reg_rdata[5] ;
 wire \u_semaphore.reg_rdata[6] ;
 wire \u_semaphore.reg_rdata[7] ;
 wire \u_semaphore.reg_rdata[8] ;
 wire \u_semaphore.reg_rdata[9] ;
 wire \u_skew_pinmux.clk_d1 ;
 wire \u_skew_pinmux.clk_d10 ;
 wire \u_skew_pinmux.clk_d11 ;
 wire \u_skew_pinmux.clk_d12 ;
 wire \u_skew_pinmux.clk_d13 ;
 wire \u_skew_pinmux.clk_d14 ;
 wire \u_skew_pinmux.clk_d15 ;
 wire \u_skew_pinmux.clk_d2 ;
 wire \u_skew_pinmux.clk_d3 ;
 wire \u_skew_pinmux.clk_d4 ;
 wire \u_skew_pinmux.clk_d5 ;
 wire \u_skew_pinmux.clk_d6 ;
 wire \u_skew_pinmux.clk_d7 ;
 wire \u_skew_pinmux.clk_d8 ;
 wire \u_skew_pinmux.clk_d9 ;
 wire \u_skew_pinmux.clk_inbuf ;
 wire \u_skew_pinmux.clkbuf_1.X1 ;
 wire \u_skew_pinmux.clkbuf_1.X2 ;
 wire \u_skew_pinmux.clkbuf_1.X3 ;
 wire \u_skew_pinmux.clkbuf_10.X1 ;
 wire \u_skew_pinmux.clkbuf_10.X2 ;
 wire \u_skew_pinmux.clkbuf_10.X3 ;
 wire \u_skew_pinmux.clkbuf_11.X1 ;
 wire \u_skew_pinmux.clkbuf_11.X2 ;
 wire \u_skew_pinmux.clkbuf_11.X3 ;
 wire \u_skew_pinmux.clkbuf_12.X1 ;
 wire \u_skew_pinmux.clkbuf_12.X2 ;
 wire \u_skew_pinmux.clkbuf_12.X3 ;
 wire \u_skew_pinmux.clkbuf_13.X1 ;
 wire \u_skew_pinmux.clkbuf_13.X2 ;
 wire \u_skew_pinmux.clkbuf_13.X3 ;
 wire \u_skew_pinmux.clkbuf_14.X1 ;
 wire \u_skew_pinmux.clkbuf_14.X2 ;
 wire \u_skew_pinmux.clkbuf_14.X3 ;
 wire \u_skew_pinmux.clkbuf_15.X1 ;
 wire \u_skew_pinmux.clkbuf_15.X2 ;
 wire \u_skew_pinmux.clkbuf_15.X3 ;
 wire \u_skew_pinmux.clkbuf_2.X1 ;
 wire \u_skew_pinmux.clkbuf_2.X2 ;
 wire \u_skew_pinmux.clkbuf_2.X3 ;
 wire \u_skew_pinmux.clkbuf_3.X1 ;
 wire \u_skew_pinmux.clkbuf_3.X2 ;
 wire \u_skew_pinmux.clkbuf_3.X3 ;
 wire \u_skew_pinmux.clkbuf_4.X1 ;
 wire \u_skew_pinmux.clkbuf_4.X2 ;
 wire \u_skew_pinmux.clkbuf_4.X3 ;
 wire \u_skew_pinmux.clkbuf_5.X1 ;
 wire \u_skew_pinmux.clkbuf_5.X2 ;
 wire \u_skew_pinmux.clkbuf_5.X3 ;
 wire \u_skew_pinmux.clkbuf_6.X1 ;
 wire \u_skew_pinmux.clkbuf_6.X2 ;
 wire \u_skew_pinmux.clkbuf_6.X3 ;
 wire \u_skew_pinmux.clkbuf_7.X1 ;
 wire \u_skew_pinmux.clkbuf_7.X2 ;
 wire \u_skew_pinmux.clkbuf_7.X3 ;
 wire \u_skew_pinmux.clkbuf_8.X1 ;
 wire \u_skew_pinmux.clkbuf_8.X2 ;
 wire \u_skew_pinmux.clkbuf_8.X3 ;
 wire \u_skew_pinmux.clkbuf_9.X1 ;
 wire \u_skew_pinmux.clkbuf_9.X2 ;
 wire \u_skew_pinmux.clkbuf_9.X3 ;
 wire \u_skew_pinmux.d00 ;
 wire \u_skew_pinmux.d01 ;
 wire \u_skew_pinmux.d02 ;
 wire \u_skew_pinmux.d03 ;
 wire \u_skew_pinmux.d04 ;
 wire \u_skew_pinmux.d05 ;
 wire \u_skew_pinmux.d06 ;
 wire \u_skew_pinmux.d07 ;
 wire \u_skew_pinmux.d10 ;
 wire \u_skew_pinmux.d11 ;
 wire \u_skew_pinmux.d12 ;
 wire \u_skew_pinmux.d13 ;
 wire \u_skew_pinmux.d20 ;
 wire \u_skew_pinmux.d21 ;
 wire \u_skew_pinmux.d30 ;
 wire \u_skew_pinmux.in0 ;
 wire \u_skew_pinmux.in1 ;
 wire \u_skew_pinmux.in10 ;
 wire \u_skew_pinmux.in11 ;
 wire \u_skew_pinmux.in12 ;
 wire \u_skew_pinmux.in13 ;
 wire \u_skew_pinmux.in14 ;
 wire \u_skew_pinmux.in15 ;
 wire \u_skew_pinmux.in2 ;
 wire \u_skew_pinmux.in3 ;
 wire \u_skew_pinmux.in4 ;
 wire \u_skew_pinmux.in5 ;
 wire \u_skew_pinmux.in6 ;
 wire \u_skew_pinmux.in7 ;
 wire \u_skew_pinmux.in8 ;
 wire \u_skew_pinmux.in9 ;
 wire \u_timer.cfg_pulse_1us[0] ;
 wire \u_timer.cfg_pulse_1us[1] ;
 wire \u_timer.cfg_pulse_1us[2] ;
 wire \u_timer.cfg_pulse_1us[3] ;
 wire \u_timer.cfg_pulse_1us[4] ;
 wire \u_timer.cfg_pulse_1us[5] ;
 wire \u_timer.cfg_pulse_1us[6] ;
 wire \u_timer.cfg_pulse_1us[7] ;
 wire \u_timer.cfg_pulse_1us[8] ;
 wire \u_timer.cfg_pulse_1us[9] ;
 wire \u_timer.cfg_timer0[0] ;
 wire \u_timer.cfg_timer0[10] ;
 wire \u_timer.cfg_timer0[11] ;
 wire \u_timer.cfg_timer0[12] ;
 wire \u_timer.cfg_timer0[13] ;
 wire \u_timer.cfg_timer0[14] ;
 wire \u_timer.cfg_timer0[15] ;
 wire \u_timer.cfg_timer0[16] ;
 wire \u_timer.cfg_timer0[17] ;
 wire \u_timer.cfg_timer0[18] ;
 wire \u_timer.cfg_timer0[1] ;
 wire \u_timer.cfg_timer0[2] ;
 wire \u_timer.cfg_timer0[3] ;
 wire \u_timer.cfg_timer0[4] ;
 wire \u_timer.cfg_timer0[5] ;
 wire \u_timer.cfg_timer0[6] ;
 wire \u_timer.cfg_timer0[7] ;
 wire \u_timer.cfg_timer0[8] ;
 wire \u_timer.cfg_timer0[9] ;
 wire \u_timer.cfg_timer1[0] ;
 wire \u_timer.cfg_timer1[10] ;
 wire \u_timer.cfg_timer1[11] ;
 wire \u_timer.cfg_timer1[12] ;
 wire \u_timer.cfg_timer1[13] ;
 wire \u_timer.cfg_timer1[14] ;
 wire \u_timer.cfg_timer1[15] ;
 wire \u_timer.cfg_timer1[16] ;
 wire \u_timer.cfg_timer1[17] ;
 wire \u_timer.cfg_timer1[18] ;
 wire \u_timer.cfg_timer1[1] ;
 wire \u_timer.cfg_timer1[2] ;
 wire \u_timer.cfg_timer1[3] ;
 wire \u_timer.cfg_timer1[4] ;
 wire \u_timer.cfg_timer1[5] ;
 wire \u_timer.cfg_timer1[6] ;
 wire \u_timer.cfg_timer1[7] ;
 wire \u_timer.cfg_timer1[8] ;
 wire \u_timer.cfg_timer1[9] ;
 wire \u_timer.cfg_timer2[0] ;
 wire \u_timer.cfg_timer2[10] ;
 wire \u_timer.cfg_timer2[11] ;
 wire \u_timer.cfg_timer2[12] ;
 wire \u_timer.cfg_timer2[13] ;
 wire \u_timer.cfg_timer2[14] ;
 wire \u_timer.cfg_timer2[15] ;
 wire \u_timer.cfg_timer2[16] ;
 wire \u_timer.cfg_timer2[17] ;
 wire \u_timer.cfg_timer2[18] ;
 wire \u_timer.cfg_timer2[1] ;
 wire \u_timer.cfg_timer2[2] ;
 wire \u_timer.cfg_timer2[3] ;
 wire \u_timer.cfg_timer2[4] ;
 wire \u_timer.cfg_timer2[5] ;
 wire \u_timer.cfg_timer2[6] ;
 wire \u_timer.cfg_timer2[7] ;
 wire \u_timer.cfg_timer2[8] ;
 wire \u_timer.cfg_timer2[9] ;
 wire \u_timer.reg_ack ;
 wire \u_timer.reg_rdata[0] ;
 wire \u_timer.reg_rdata[10] ;
 wire \u_timer.reg_rdata[11] ;
 wire \u_timer.reg_rdata[12] ;
 wire \u_timer.reg_rdata[13] ;
 wire \u_timer.reg_rdata[14] ;
 wire \u_timer.reg_rdata[15] ;
 wire \u_timer.reg_rdata[16] ;
 wire \u_timer.reg_rdata[17] ;
 wire \u_timer.reg_rdata[18] ;
 wire \u_timer.reg_rdata[19] ;
 wire \u_timer.reg_rdata[1] ;
 wire \u_timer.reg_rdata[20] ;
 wire \u_timer.reg_rdata[21] ;
 wire \u_timer.reg_rdata[22] ;
 wire \u_timer.reg_rdata[23] ;
 wire \u_timer.reg_rdata[24] ;
 wire \u_timer.reg_rdata[25] ;
 wire \u_timer.reg_rdata[26] ;
 wire \u_timer.reg_rdata[27] ;
 wire \u_timer.reg_rdata[28] ;
 wire \u_timer.reg_rdata[29] ;
 wire \u_timer.reg_rdata[2] ;
 wire \u_timer.reg_rdata[30] ;
 wire \u_timer.reg_rdata[31] ;
 wire \u_timer.reg_rdata[3] ;
 wire \u_timer.reg_rdata[4] ;
 wire \u_timer.reg_rdata[5] ;
 wire \u_timer.reg_rdata[6] ;
 wire \u_timer.reg_rdata[7] ;
 wire \u_timer.reg_rdata[8] ;
 wire \u_timer.reg_rdata[9] ;
 wire \u_timer.u_pulse_1ms.cnt[0] ;
 wire \u_timer.u_pulse_1ms.cnt[1] ;
 wire \u_timer.u_pulse_1ms.cnt[2] ;
 wire \u_timer.u_pulse_1ms.cnt[3] ;
 wire \u_timer.u_pulse_1ms.cnt[4] ;
 wire \u_timer.u_pulse_1ms.cnt[5] ;
 wire \u_timer.u_pulse_1ms.cnt[6] ;
 wire \u_timer.u_pulse_1ms.cnt[7] ;
 wire \u_timer.u_pulse_1ms.cnt[8] ;
 wire \u_timer.u_pulse_1ms.cnt[9] ;
 wire \u_timer.u_pulse_1s.cnt[0] ;
 wire \u_timer.u_pulse_1s.cnt[1] ;
 wire \u_timer.u_pulse_1s.cnt[2] ;
 wire \u_timer.u_pulse_1s.cnt[3] ;
 wire \u_timer.u_pulse_1s.cnt[4] ;
 wire \u_timer.u_pulse_1s.cnt[5] ;
 wire \u_timer.u_pulse_1s.cnt[6] ;
 wire \u_timer.u_pulse_1s.cnt[7] ;
 wire \u_timer.u_pulse_1s.cnt[8] ;
 wire \u_timer.u_pulse_1s.cnt[9] ;
 wire \u_timer.u_pulse_1us.cnt[0] ;
 wire \u_timer.u_pulse_1us.cnt[1] ;
 wire \u_timer.u_pulse_1us.cnt[2] ;
 wire \u_timer.u_pulse_1us.cnt[3] ;
 wire \u_timer.u_pulse_1us.cnt[4] ;
 wire \u_timer.u_pulse_1us.cnt[5] ;
 wire \u_timer.u_pulse_1us.cnt[6] ;
 wire \u_timer.u_pulse_1us.cnt[7] ;
 wire \u_timer.u_pulse_1us.cnt[8] ;
 wire \u_timer.u_pulse_1us.cnt[9] ;
 wire \u_timer.u_reg.reg_0[10] ;
 wire \u_timer.u_reg.reg_0[11] ;
 wire \u_timer.u_reg.reg_0[12] ;
 wire \u_timer.u_reg.reg_0[13] ;
 wire \u_timer.u_reg.reg_0[14] ;
 wire \u_timer.u_reg.reg_0[15] ;
 wire \u_timer.u_reg.reg_0[16] ;
 wire \u_timer.u_reg.reg_0[17] ;
 wire \u_timer.u_reg.reg_0[18] ;
 wire \u_timer.u_reg.reg_0[19] ;
 wire \u_timer.u_reg.reg_0[20] ;
 wire \u_timer.u_reg.reg_0[21] ;
 wire \u_timer.u_reg.reg_0[22] ;
 wire \u_timer.u_reg.reg_0[23] ;
 wire \u_timer.u_reg.reg_0[24] ;
 wire \u_timer.u_reg.reg_0[25] ;
 wire \u_timer.u_reg.reg_0[26] ;
 wire \u_timer.u_reg.reg_0[27] ;
 wire \u_timer.u_reg.reg_0[28] ;
 wire \u_timer.u_reg.reg_0[29] ;
 wire \u_timer.u_reg.reg_0[30] ;
 wire \u_timer.u_reg.reg_0[31] ;
 wire \u_timer.u_reg.reg_1[19] ;
 wire \u_timer.u_reg.reg_1[20] ;
 wire \u_timer.u_reg.reg_1[21] ;
 wire \u_timer.u_reg.reg_1[22] ;
 wire \u_timer.u_reg.reg_1[23] ;
 wire \u_timer.u_reg.reg_1[24] ;
 wire \u_timer.u_reg.reg_1[25] ;
 wire \u_timer.u_reg.reg_1[26] ;
 wire \u_timer.u_reg.reg_1[27] ;
 wire \u_timer.u_reg.reg_1[28] ;
 wire \u_timer.u_reg.reg_1[29] ;
 wire \u_timer.u_reg.reg_1[30] ;
 wire \u_timer.u_reg.reg_1[31] ;
 wire \u_timer.u_reg.reg_2[19] ;
 wire \u_timer.u_reg.reg_2[20] ;
 wire \u_timer.u_reg.reg_2[21] ;
 wire \u_timer.u_reg.reg_2[22] ;
 wire \u_timer.u_reg.reg_2[23] ;
 wire \u_timer.u_reg.reg_2[24] ;
 wire \u_timer.u_reg.reg_2[25] ;
 wire \u_timer.u_reg.reg_2[26] ;
 wire \u_timer.u_reg.reg_2[27] ;
 wire \u_timer.u_reg.reg_2[28] ;
 wire \u_timer.u_reg.reg_2[29] ;
 wire \u_timer.u_reg.reg_2[30] ;
 wire \u_timer.u_reg.reg_2[31] ;
 wire \u_timer.u_reg.reg_3[19] ;
 wire \u_timer.u_reg.reg_3[20] ;
 wire \u_timer.u_reg.reg_3[21] ;
 wire \u_timer.u_reg.reg_3[22] ;
 wire \u_timer.u_reg.reg_3[23] ;
 wire \u_timer.u_reg.reg_3[24] ;
 wire \u_timer.u_reg.reg_3[25] ;
 wire \u_timer.u_reg.reg_3[26] ;
 wire \u_timer.u_reg.reg_3[27] ;
 wire \u_timer.u_reg.reg_3[28] ;
 wire \u_timer.u_reg.reg_3[29] ;
 wire \u_timer.u_reg.reg_3[30] ;
 wire \u_timer.u_reg.reg_3[31] ;
 wire \u_timer.u_reg.reg_out[0] ;
 wire \u_timer.u_reg.reg_out[10] ;
 wire \u_timer.u_reg.reg_out[11] ;
 wire \u_timer.u_reg.reg_out[12] ;
 wire \u_timer.u_reg.reg_out[13] ;
 wire \u_timer.u_reg.reg_out[14] ;
 wire \u_timer.u_reg.reg_out[15] ;
 wire \u_timer.u_reg.reg_out[16] ;
 wire \u_timer.u_reg.reg_out[17] ;
 wire \u_timer.u_reg.reg_out[18] ;
 wire \u_timer.u_reg.reg_out[19] ;
 wire \u_timer.u_reg.reg_out[1] ;
 wire \u_timer.u_reg.reg_out[20] ;
 wire \u_timer.u_reg.reg_out[21] ;
 wire \u_timer.u_reg.reg_out[22] ;
 wire \u_timer.u_reg.reg_out[23] ;
 wire \u_timer.u_reg.reg_out[24] ;
 wire \u_timer.u_reg.reg_out[25] ;
 wire \u_timer.u_reg.reg_out[26] ;
 wire \u_timer.u_reg.reg_out[27] ;
 wire \u_timer.u_reg.reg_out[28] ;
 wire \u_timer.u_reg.reg_out[29] ;
 wire \u_timer.u_reg.reg_out[2] ;
 wire \u_timer.u_reg.reg_out[30] ;
 wire \u_timer.u_reg.reg_out[31] ;
 wire \u_timer.u_reg.reg_out[3] ;
 wire \u_timer.u_reg.reg_out[4] ;
 wire \u_timer.u_reg.reg_out[5] ;
 wire \u_timer.u_reg.reg_out[6] ;
 wire \u_timer.u_reg.reg_out[7] ;
 wire \u_timer.u_reg.reg_out[8] ;
 wire \u_timer.u_reg.reg_out[9] ;
 wire \u_timer.u_timer_0.timer_counter[0] ;
 wire \u_timer.u_timer_0.timer_counter[10] ;
 wire \u_timer.u_timer_0.timer_counter[11] ;
 wire \u_timer.u_timer_0.timer_counter[12] ;
 wire \u_timer.u_timer_0.timer_counter[13] ;
 wire \u_timer.u_timer_0.timer_counter[14] ;
 wire \u_timer.u_timer_0.timer_counter[15] ;
 wire \u_timer.u_timer_0.timer_counter[1] ;
 wire \u_timer.u_timer_0.timer_counter[2] ;
 wire \u_timer.u_timer_0.timer_counter[3] ;
 wire \u_timer.u_timer_0.timer_counter[4] ;
 wire \u_timer.u_timer_0.timer_counter[5] ;
 wire \u_timer.u_timer_0.timer_counter[6] ;
 wire \u_timer.u_timer_0.timer_counter[7] ;
 wire \u_timer.u_timer_0.timer_counter[8] ;
 wire \u_timer.u_timer_0.timer_counter[9] ;
 wire \u_timer.u_timer_0.timer_hit ;
 wire \u_timer.u_timer_0.timer_hit_s1 ;
 wire \u_timer.u_timer_1.timer_counter[0] ;
 wire \u_timer.u_timer_1.timer_counter[10] ;
 wire \u_timer.u_timer_1.timer_counter[11] ;
 wire \u_timer.u_timer_1.timer_counter[12] ;
 wire \u_timer.u_timer_1.timer_counter[13] ;
 wire \u_timer.u_timer_1.timer_counter[14] ;
 wire \u_timer.u_timer_1.timer_counter[15] ;
 wire \u_timer.u_timer_1.timer_counter[1] ;
 wire \u_timer.u_timer_1.timer_counter[2] ;
 wire \u_timer.u_timer_1.timer_counter[3] ;
 wire \u_timer.u_timer_1.timer_counter[4] ;
 wire \u_timer.u_timer_1.timer_counter[5] ;
 wire \u_timer.u_timer_1.timer_counter[6] ;
 wire \u_timer.u_timer_1.timer_counter[7] ;
 wire \u_timer.u_timer_1.timer_counter[8] ;
 wire \u_timer.u_timer_1.timer_counter[9] ;
 wire \u_timer.u_timer_1.timer_hit ;
 wire \u_timer.u_timer_1.timer_hit_s1 ;
 wire \u_timer.u_timer_2.timer_counter[0] ;
 wire \u_timer.u_timer_2.timer_counter[10] ;
 wire \u_timer.u_timer_2.timer_counter[11] ;
 wire \u_timer.u_timer_2.timer_counter[12] ;
 wire \u_timer.u_timer_2.timer_counter[13] ;
 wire \u_timer.u_timer_2.timer_counter[14] ;
 wire \u_timer.u_timer_2.timer_counter[15] ;
 wire \u_timer.u_timer_2.timer_counter[1] ;
 wire \u_timer.u_timer_2.timer_counter[2] ;
 wire \u_timer.u_timer_2.timer_counter[3] ;
 wire \u_timer.u_timer_2.timer_counter[4] ;
 wire \u_timer.u_timer_2.timer_counter[5] ;
 wire \u_timer.u_timer_2.timer_counter[6] ;
 wire \u_timer.u_timer_2.timer_counter[7] ;
 wire \u_timer.u_timer_2.timer_counter[8] ;
 wire \u_timer.u_timer_2.timer_counter[9] ;
 wire \u_timer.u_timer_2.timer_hit ;
 wire \u_timer.u_timer_2.timer_hit_s1 ;
 wire \u_ws281x.cfg_clk_period[0] ;
 wire \u_ws281x.cfg_clk_period[1] ;
 wire \u_ws281x.cfg_clk_period[2] ;
 wire \u_ws281x.cfg_clk_period[3] ;
 wire \u_ws281x.cfg_clk_period[4] ;
 wire \u_ws281x.cfg_clk_period[5] ;
 wire \u_ws281x.cfg_clk_period[6] ;
 wire \u_ws281x.cfg_clk_period[7] ;
 wire \u_ws281x.cfg_clk_period[8] ;
 wire \u_ws281x.cfg_clk_period[9] ;
 wire \u_ws281x.cfg_reset_period[0] ;
 wire \u_ws281x.cfg_reset_period[10] ;
 wire \u_ws281x.cfg_reset_period[11] ;
 wire \u_ws281x.cfg_reset_period[12] ;
 wire \u_ws281x.cfg_reset_period[13] ;
 wire \u_ws281x.cfg_reset_period[14] ;
 wire \u_ws281x.cfg_reset_period[15] ;
 wire \u_ws281x.cfg_reset_period[1] ;
 wire \u_ws281x.cfg_reset_period[2] ;
 wire \u_ws281x.cfg_reset_period[3] ;
 wire \u_ws281x.cfg_reset_period[4] ;
 wire \u_ws281x.cfg_reset_period[5] ;
 wire \u_ws281x.cfg_reset_period[6] ;
 wire \u_ws281x.cfg_reset_period[7] ;
 wire \u_ws281x.cfg_reset_period[8] ;
 wire \u_ws281x.cfg_reset_period[9] ;
 wire \u_ws281x.cfg_th0_period[0] ;
 wire \u_ws281x.cfg_th0_period[1] ;
 wire \u_ws281x.cfg_th0_period[2] ;
 wire \u_ws281x.cfg_th0_period[3] ;
 wire \u_ws281x.cfg_th0_period[4] ;
 wire \u_ws281x.cfg_th0_period[5] ;
 wire \u_ws281x.cfg_th0_period[6] ;
 wire \u_ws281x.cfg_th0_period[7] ;
 wire \u_ws281x.cfg_th0_period[8] ;
 wire \u_ws281x.cfg_th0_period[9] ;
 wire \u_ws281x.cfg_th1_period[0] ;
 wire \u_ws281x.cfg_th1_period[1] ;
 wire \u_ws281x.cfg_th1_period[2] ;
 wire \u_ws281x.cfg_th1_period[3] ;
 wire \u_ws281x.cfg_th1_period[4] ;
 wire \u_ws281x.cfg_th1_period[5] ;
 wire \u_ws281x.cfg_th1_period[6] ;
 wire \u_ws281x.cfg_th1_period[7] ;
 wire \u_ws281x.cfg_th1_period[8] ;
 wire \u_ws281x.cfg_th1_period[9] ;
 wire \u_ws281x.port0_enb ;
 wire \u_ws281x.port0_rd ;
 wire \u_ws281x.port1_enb ;
 wire \u_ws281x.port1_rd ;
 wire \u_ws281x.reg_ack ;
 wire \u_ws281x.reg_rdata[0] ;
 wire \u_ws281x.reg_rdata[10] ;
 wire \u_ws281x.reg_rdata[11] ;
 wire \u_ws281x.reg_rdata[12] ;
 wire \u_ws281x.reg_rdata[13] ;
 wire \u_ws281x.reg_rdata[14] ;
 wire \u_ws281x.reg_rdata[15] ;
 wire \u_ws281x.reg_rdata[16] ;
 wire \u_ws281x.reg_rdata[17] ;
 wire \u_ws281x.reg_rdata[18] ;
 wire \u_ws281x.reg_rdata[19] ;
 wire \u_ws281x.reg_rdata[1] ;
 wire \u_ws281x.reg_rdata[20] ;
 wire \u_ws281x.reg_rdata[21] ;
 wire \u_ws281x.reg_rdata[22] ;
 wire \u_ws281x.reg_rdata[23] ;
 wire \u_ws281x.reg_rdata[24] ;
 wire \u_ws281x.reg_rdata[25] ;
 wire \u_ws281x.reg_rdata[26] ;
 wire \u_ws281x.reg_rdata[27] ;
 wire \u_ws281x.reg_rdata[28] ;
 wire \u_ws281x.reg_rdata[29] ;
 wire \u_ws281x.reg_rdata[2] ;
 wire \u_ws281x.reg_rdata[30] ;
 wire \u_ws281x.reg_rdata[31] ;
 wire \u_ws281x.reg_rdata[3] ;
 wire \u_ws281x.reg_rdata[4] ;
 wire \u_ws281x.reg_rdata[5] ;
 wire \u_ws281x.reg_rdata[6] ;
 wire \u_ws281x.reg_rdata[7] ;
 wire \u_ws281x.reg_rdata[8] ;
 wire \u_ws281x.reg_rdata[9] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.empty ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.full ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][0] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][10] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][11] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][12] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][13] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][14] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][15] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][16] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][17] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][18] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][19] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][1] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][20] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][21] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][22] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][23] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][2] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][3] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][4] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][5] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][6] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][7] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][8] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][9] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][0] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][10] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][11] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][12] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][13] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][14] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][15] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][16] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][17] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][18] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][19] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][1] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][20] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][21] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][22] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][23] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][2] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][3] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][4] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][5] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][6] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][7] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][8] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][9] ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.rd_ptr ;
 wire \u_ws281x.u_reg.gfifo[0].u_fifo.wr_ptr ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.empty ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.full ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][0] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][10] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][11] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][12] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][13] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][14] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][15] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][16] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][17] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][18] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][19] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][1] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][20] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][21] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][22] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][23] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][2] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][3] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][4] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][5] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][6] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][7] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][8] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][9] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][0] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][10] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][11] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][12] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][13] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][14] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][15] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][16] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][17] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][18] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][19] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][1] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][20] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][21] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][22] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][23] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][2] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][3] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][4] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][5] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][6] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][7] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][8] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][9] ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.rd_ptr ;
 wire \u_ws281x.u_reg.gfifo[1].u_fifo.wr_ptr ;
 wire \u_ws281x.u_reg.reg_2[30] ;
 wire \u_ws281x.u_reg.reg_2[31] ;
 wire \u_ws281x.u_reg.reg_out[0] ;
 wire \u_ws281x.u_reg.reg_out[10] ;
 wire \u_ws281x.u_reg.reg_out[11] ;
 wire \u_ws281x.u_reg.reg_out[12] ;
 wire \u_ws281x.u_reg.reg_out[13] ;
 wire \u_ws281x.u_reg.reg_out[14] ;
 wire \u_ws281x.u_reg.reg_out[15] ;
 wire \u_ws281x.u_reg.reg_out[16] ;
 wire \u_ws281x.u_reg.reg_out[17] ;
 wire \u_ws281x.u_reg.reg_out[18] ;
 wire \u_ws281x.u_reg.reg_out[19] ;
 wire \u_ws281x.u_reg.reg_out[1] ;
 wire \u_ws281x.u_reg.reg_out[20] ;
 wire \u_ws281x.u_reg.reg_out[21] ;
 wire \u_ws281x.u_reg.reg_out[22] ;
 wire \u_ws281x.u_reg.reg_out[23] ;
 wire \u_ws281x.u_reg.reg_out[24] ;
 wire \u_ws281x.u_reg.reg_out[25] ;
 wire \u_ws281x.u_reg.reg_out[26] ;
 wire \u_ws281x.u_reg.reg_out[27] ;
 wire \u_ws281x.u_reg.reg_out[28] ;
 wire \u_ws281x.u_reg.reg_out[29] ;
 wire \u_ws281x.u_reg.reg_out[2] ;
 wire \u_ws281x.u_reg.reg_out[30] ;
 wire \u_ws281x.u_reg.reg_out[31] ;
 wire \u_ws281x.u_reg.reg_out[3] ;
 wire \u_ws281x.u_reg.reg_out[4] ;
 wire \u_ws281x.u_reg.reg_out[5] ;
 wire \u_ws281x.u_reg.reg_out[6] ;
 wire \u_ws281x.u_reg.reg_out[7] ;
 wire \u_ws281x.u_reg.reg_out[8] ;
 wire \u_ws281x.u_reg.reg_out[9] ;
 wire \u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ;
 wire \u_ws281x.u_reg.u_reg_0.gen_bit_reg[2].u_bit_reg.data_out ;
 wire \u_ws281x.u_reg.u_reg_0.gen_bit_reg[3].u_bit_reg.data_out ;
 wire \u_ws281x.u_txd_0.bit_cnt[0] ;
 wire \u_ws281x.u_txd_0.bit_cnt[1] ;
 wire \u_ws281x.u_txd_0.bit_cnt[2] ;
 wire \u_ws281x.u_txd_0.bit_cnt[3] ;
 wire \u_ws281x.u_txd_0.bit_cnt[4] ;
 wire \u_ws281x.u_txd_0.clk_cnt[0] ;
 wire \u_ws281x.u_txd_0.clk_cnt[10] ;
 wire \u_ws281x.u_txd_0.clk_cnt[11] ;
 wire \u_ws281x.u_txd_0.clk_cnt[12] ;
 wire \u_ws281x.u_txd_0.clk_cnt[13] ;
 wire \u_ws281x.u_txd_0.clk_cnt[14] ;
 wire \u_ws281x.u_txd_0.clk_cnt[15] ;
 wire \u_ws281x.u_txd_0.clk_cnt[1] ;
 wire \u_ws281x.u_txd_0.clk_cnt[2] ;
 wire \u_ws281x.u_txd_0.clk_cnt[3] ;
 wire \u_ws281x.u_txd_0.clk_cnt[4] ;
 wire \u_ws281x.u_txd_0.clk_cnt[5] ;
 wire \u_ws281x.u_txd_0.clk_cnt[6] ;
 wire \u_ws281x.u_txd_0.clk_cnt[7] ;
 wire \u_ws281x.u_txd_0.clk_cnt[8] ;
 wire \u_ws281x.u_txd_0.clk_cnt[9] ;
 wire \u_ws281x.u_txd_0.led_data[0] ;
 wire \u_ws281x.u_txd_0.led_data[10] ;
 wire \u_ws281x.u_txd_0.led_data[11] ;
 wire \u_ws281x.u_txd_0.led_data[12] ;
 wire \u_ws281x.u_txd_0.led_data[13] ;
 wire \u_ws281x.u_txd_0.led_data[14] ;
 wire \u_ws281x.u_txd_0.led_data[15] ;
 wire \u_ws281x.u_txd_0.led_data[16] ;
 wire \u_ws281x.u_txd_0.led_data[17] ;
 wire \u_ws281x.u_txd_0.led_data[18] ;
 wire \u_ws281x.u_txd_0.led_data[19] ;
 wire \u_ws281x.u_txd_0.led_data[1] ;
 wire \u_ws281x.u_txd_0.led_data[20] ;
 wire \u_ws281x.u_txd_0.led_data[21] ;
 wire \u_ws281x.u_txd_0.led_data[22] ;
 wire \u_ws281x.u_txd_0.led_data[23] ;
 wire \u_ws281x.u_txd_0.led_data[2] ;
 wire \u_ws281x.u_txd_0.led_data[3] ;
 wire \u_ws281x.u_txd_0.led_data[4] ;
 wire \u_ws281x.u_txd_0.led_data[5] ;
 wire \u_ws281x.u_txd_0.led_data[6] ;
 wire \u_ws281x.u_txd_0.led_data[7] ;
 wire \u_ws281x.u_txd_0.led_data[8] ;
 wire \u_ws281x.u_txd_0.led_data[9] ;
 wire \u_ws281x.u_txd_0.state ;
 wire \u_ws281x.u_txd_0.txd ;
 wire \u_ws281x.u_txd_1.bit_cnt[0] ;
 wire \u_ws281x.u_txd_1.bit_cnt[1] ;
 wire \u_ws281x.u_txd_1.bit_cnt[2] ;
 wire \u_ws281x.u_txd_1.bit_cnt[3] ;
 wire \u_ws281x.u_txd_1.bit_cnt[4] ;
 wire \u_ws281x.u_txd_1.clk_cnt[0] ;
 wire \u_ws281x.u_txd_1.clk_cnt[10] ;
 wire \u_ws281x.u_txd_1.clk_cnt[11] ;
 wire \u_ws281x.u_txd_1.clk_cnt[12] ;
 wire \u_ws281x.u_txd_1.clk_cnt[13] ;
 wire \u_ws281x.u_txd_1.clk_cnt[14] ;
 wire \u_ws281x.u_txd_1.clk_cnt[15] ;
 wire \u_ws281x.u_txd_1.clk_cnt[1] ;
 wire \u_ws281x.u_txd_1.clk_cnt[2] ;
 wire \u_ws281x.u_txd_1.clk_cnt[3] ;
 wire \u_ws281x.u_txd_1.clk_cnt[4] ;
 wire \u_ws281x.u_txd_1.clk_cnt[5] ;
 wire \u_ws281x.u_txd_1.clk_cnt[6] ;
 wire \u_ws281x.u_txd_1.clk_cnt[7] ;
 wire \u_ws281x.u_txd_1.clk_cnt[8] ;
 wire \u_ws281x.u_txd_1.clk_cnt[9] ;
 wire \u_ws281x.u_txd_1.led_data[0] ;
 wire \u_ws281x.u_txd_1.led_data[10] ;
 wire \u_ws281x.u_txd_1.led_data[11] ;
 wire \u_ws281x.u_txd_1.led_data[12] ;
 wire \u_ws281x.u_txd_1.led_data[13] ;
 wire \u_ws281x.u_txd_1.led_data[14] ;
 wire \u_ws281x.u_txd_1.led_data[15] ;
 wire \u_ws281x.u_txd_1.led_data[16] ;
 wire \u_ws281x.u_txd_1.led_data[17] ;
 wire \u_ws281x.u_txd_1.led_data[18] ;
 wire \u_ws281x.u_txd_1.led_data[19] ;
 wire \u_ws281x.u_txd_1.led_data[1] ;
 wire \u_ws281x.u_txd_1.led_data[20] ;
 wire \u_ws281x.u_txd_1.led_data[21] ;
 wire \u_ws281x.u_txd_1.led_data[22] ;
 wire \u_ws281x.u_txd_1.led_data[23] ;
 wire \u_ws281x.u_txd_1.led_data[2] ;
 wire \u_ws281x.u_txd_1.led_data[3] ;
 wire \u_ws281x.u_txd_1.led_data[4] ;
 wire \u_ws281x.u_txd_1.led_data[5] ;
 wire \u_ws281x.u_txd_1.led_data[6] ;
 wire \u_ws281x.u_txd_1.led_data[7] ;
 wire \u_ws281x.u_txd_1.led_data[8] ;
 wire \u_ws281x.u_txd_1.led_data[9] ;
 wire \u_ws281x.u_txd_1.state ;
 wire \u_ws281x.u_txd_1.txd ;

 sky130_fd_sc_hd__diode_2 ANTENNA__04690__A (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__04691__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__04692__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__04693__A (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__04694__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__04701__A (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04702__A (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04704__A (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04710__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__04711__A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__04715__A (.DIODE(\u_ws281x.cfg_clk_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04717__A (.DIODE(\u_ws281x.cfg_clk_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04722__A (.DIODE(\u_ws281x.cfg_clk_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04725__A (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04728__A (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04729__A (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04730__A (.DIODE(\u_ws281x.cfg_reset_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04731__A (.DIODE(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04733__A (.DIODE(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04736__A (.DIODE(\u_ws281x.cfg_reset_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04740__A (.DIODE(\u_ws281x.cfg_reset_period[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04749__A (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04751__A (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04753__A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04754__A (.DIODE(\u_ws281x.port1_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04766__A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.full ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04768__A (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__04770__A (.DIODE(\u_ws281x.cfg_th0_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04772__A (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04775__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__04776__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04777__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04778__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04779__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04781__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04787__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04796__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04797__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04799__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04800__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04801__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04802__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04804__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04806__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04807__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04809__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04810__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04817__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04818__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04821__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04857__A (.DIODE(\u_gpio.cfg_gpio_dir_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04858__A (.DIODE(\u_gpio.cfg_gpio_dir_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04861__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04871__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04872__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04885__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04898__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04904__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__04906__A (.DIODE(net1651));
 sky130_fd_sc_hd__diode_2 ANTENNA__04907__A (.DIODE(net1403));
 sky130_fd_sc_hd__diode_2 ANTENNA__04910__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04911__B (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04912__B1 (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04914__A_N (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04915__A (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04916__S (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04917__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04917__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__04918__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04918__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__04919__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__04919__B (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__04920__A (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__04920__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__04921__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__04922__B (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04923__A_N (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__04923__B (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__04924__A (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__04924__B (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__B (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__C (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04925__D (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04926__A (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04926__B (.DIODE(_01001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04926__C (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__04927__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__04927__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04928__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__04928__B (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__04929__A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__04929__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__04930__B (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__A1 (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__A2 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__A3 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__A4 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__04931__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04932__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__04932__A2 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04936__B1 (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__04936__B2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__A (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__B (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__C (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__04938__D (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__04939__A1 (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__04939__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04943__B2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__04945__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04949__B1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__04949__B2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__04951__A1 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__04951__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04955__B1 (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__04955__B2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04957__A1 (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__04957__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04961__B1 (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__04961__B2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04963__A1 (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__04963__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04967__B1 (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__04967__B2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04969__A1 (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__04969__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04970__B1 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04972__A_N (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04972__C (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04973__A3 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04974__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__04974__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__A1 (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__A2 (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__A3 (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__A4 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__04975__B1 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__04976__A1 (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__04976__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__04977__B1 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04979__A_N (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04979__C (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04980__A3 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04981__A1 (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__04981__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__04982__A1 (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__04982__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__04985__A_N (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04986__A3 (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__04987__A1 (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__04987__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__04988__A1 (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__04988__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__04991__A (.DIODE(_01040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04993__A3 (.DIODE(_01040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__04994__A1 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__04994__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__04995__A1 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__04995__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__05001__A1 (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05001__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__05002__A1 (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05002__A2 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05003__B1 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05005__A_N (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05005__C (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05006__A3 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05007__A1 (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__05007__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__05008__A1 (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__05008__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__05011__A_N (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05012__A3 (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05013__A1 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__05013__A2 (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__05014__A1 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__05014__A2 (.DIODE(net535));
 sky130_fd_sc_hd__diode_2 ANTENNA__05017__A_N (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05018__A3 (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05019__A1 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__05019__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05020__A1 (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__05020__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05021__A (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__05021__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__05022__A (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__05022__B (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05023__B1 (.DIODE(\u_gpio.u_bit[24].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05025__A_N (.DIODE(\u_gpio.u_bit[24].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05026__A (.DIODE(\u_gpio.u_bit[24].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05028__A1 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__05028__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05029__A1 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__05029__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05030__B1 (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05032__A_N (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05033__A (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05034__S (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05035__A1 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__05035__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05036__A1 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__05036__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05037__B1 (.DIODE(\u_gpio.u_bit[26].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05039__A_N (.DIODE(\u_gpio.u_bit[26].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05040__A (.DIODE(\u_gpio.u_bit[26].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05042__A1 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__05042__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05043__A1 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__05043__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05044__B1 (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05046__A_N (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05047__A (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05048__S (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05049__A1 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__05049__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05050__A1 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__05050__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05051__B1 (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05053__A_N (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05054__A (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05055__S (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05056__A1 (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__05056__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05057__A1 (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__05057__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05058__B1 (.DIODE(\u_gpio.u_bit[29].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05060__A_N (.DIODE(\u_gpio.u_bit[29].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05061__A (.DIODE(\u_gpio.u_bit[29].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05063__A1 (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__05063__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A1 (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__05064__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05070__A1 (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__05070__A2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05071__A1 (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__05071__A2 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05077__A1 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__05077__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05078__A1 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__05078__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05079__B1 (.DIODE(\u_gpio.u_bit[31].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05081__A_N (.DIODE(\u_gpio.u_bit[31].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05082__A (.DIODE(\u_gpio.u_bit[31].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05084__A1 (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__05084__A2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05085__A1 (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__05085__A2 (.DIODE(net534));
 sky130_fd_sc_hd__diode_2 ANTENNA__05091__A1 (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__05091__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__05092__A1 (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__05092__A2 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05093__B1 (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05095__A_N (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05096__A (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05097__S (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05098__A1 (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__05098__A2 (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__05099__A1 (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__05099__A2 (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05100__A (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__05100__B (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05101__A (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__05101__B (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05102__A (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__05102__B (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA__05103__A (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__05103__B (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05104__A (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__05104__B (.DIODE(net576));
 sky130_fd_sc_hd__diode_2 ANTENNA__05105__A (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__05105__B (.DIODE(_01009_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05109__B2 (.DIODE(net577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05111__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05115__B1 (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__05115__B2 (.DIODE(net575));
 sky130_fd_sc_hd__diode_2 ANTENNA__05117__A1 (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__05117__A2 (.DIODE(_01013_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05129__A_N (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05129__B (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05129__C (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05129__D (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__05130__A (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__05130__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__05131__A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__05131__B (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__05132__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05132__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__05133__A (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05133__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__05134__A (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__05135__A (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05135__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05135__C (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__05135__D (.DIODE(_01118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05136__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05136__B (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05137__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05137__B2 (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__05138__A (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05138__C (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__05138__D (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05139__A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__05139__B (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05140__A1 (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__05140__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05141__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05142__A1 (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__05142__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05143__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05143__B (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05144__A1 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05144__A2 (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA__05144__A3 (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05144__B1 (.DIODE(\u_glbl_reg.ir_intr_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05145__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__05145__B (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05146__A1 (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA__05146__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05147__A1 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05147__A2 (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__05147__A3 (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05147__B1 (.DIODE(\u_glbl_reg.rtc_intr_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05148__A1 (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA__05148__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05149__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05149__B (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05150__B2 (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__05151__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05151__B (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05152__A1 (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__05153__B2 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__05154__A1 (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__05155__B2 (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__05156__A1 (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__05157__B2 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__05158__A1 (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__05159__B2 (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__05160__A1 (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__05161__B2 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__05162__A1 (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__05163__B2 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__05164__A1 (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__05165__B2 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__05166__A1 (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__05167__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05167__B (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05168__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05168__B2 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__05169__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05169__B (.DIODE(_01121_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05170__A1 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__05171__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05172__A1 (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__05173__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05173__B2 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__05174__A1 (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__05175__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05175__B2 (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__05177__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05177__B2 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__05178__A1 (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__05179__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05179__B2 (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__05180__A1 (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__05181__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05181__B2 (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__05182__A1 (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__05183__B1 (.DIODE(_01127_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05183__B2 (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__05184__A1 (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__05185__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05185__B2 (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__05186__A1 (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__05186__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05187__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05187__B2 (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__05188__A1 (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__05188__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05189__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05190__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05191__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05191__B2 (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__05192__A1 (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__05192__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05193__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05194__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05195__B1 (.DIODE(_01120_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05195__B2 (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__05196__A1 (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__05196__A2 (.DIODE(_01122_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05197__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__05197__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__05198__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__05198__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__05199__A (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05200__B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__05200__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05201__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05201__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05201__A3 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__05202__A1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05202__A2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05202__A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__05202__B1 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__A1 (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__A2 (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__A3 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__05203__B1 (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05204__A1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05204__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05204__A3 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__05205__A (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05206__B (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__05206__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05207__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05207__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05207__A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__05207__B1 (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__A1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__A2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__A3 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__05208__B1 (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05209__A1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05209__A2 (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05209__A3 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__05209__B1 (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__A1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__A2 (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__A3 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__05210__B1 (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05222__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__05222__B (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__05223__A (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA__05223__B (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05224__A (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05224__B (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__A2 (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__A3 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__B1 (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05225__C1 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05226__A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__05226__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05226__C (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__05227__A1 (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05227__A2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05227__B1 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05228__A1 (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05228__A2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05228__B1 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05229__A1 (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05229__A2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05229__B1 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05230__A1 (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05230__A2 (.DIODE(_01147_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05230__B1 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05243__B1 (.DIODE(_00821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05243__B2 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05244__A1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05245__A2 (.DIODE(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05245__B1 (.DIODE(_00821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05245__B2 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05246__A2 (.DIODE(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05246__B1 (.DIODE(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05248__A2_N (.DIODE(_00822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05249__B (.DIODE(\u_ws281x.cfg_reset_period[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05250__A2 (.DIODE(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05251__A1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05252__B (.DIODE(\u_ws281x.cfg_reset_period[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__A2 (.DIODE(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05253__B1 (.DIODE(\u_ws281x.cfg_reset_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05254__A2 (.DIODE(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05255__A2 (.DIODE(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05255__B1 (.DIODE(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05257__B2 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05258__A2 (.DIODE(_00822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05259__A2 (.DIODE(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05260__A2 (.DIODE(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05265__A1 (.DIODE(\u_ws281x.cfg_clk_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05265__B2 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05266__A1_N (.DIODE(\u_ws281x.cfg_clk_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05268__B1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05272__B1 (.DIODE(\u_ws281x.cfg_clk_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05273__A1 (.DIODE(\u_ws281x.cfg_clk_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05284__A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__05285__A1 (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05285__C1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__05286__A (.DIODE(\u_ws281x.cfg_reset_period[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05287__A1 (.DIODE(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05288__A1 (.DIODE(\u_ws281x.cfg_reset_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05288__B2 (.DIODE(_00822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05289__A1 (.DIODE(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05289__B2 (.DIODE(_00821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05290__A1 (.DIODE(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05290__B2 (.DIODE(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05291__B2 (.DIODE(_00821_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05293__A2 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05295__A (.DIODE(\u_ws281x.cfg_reset_period[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05296__B1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05297__A1 (.DIODE(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05298__A1 (.DIODE(\u_ws281x.cfg_reset_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05299__A1 (.DIODE(_00822_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05300__A1 (.DIODE(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05301__A1 (.DIODE(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05302__A1 (.DIODE(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05306__A (.DIODE(\u_ws281x.port1_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05310__A1 (.DIODE(\u_ws281x.cfg_clk_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05312__A (.DIODE(\u_ws281x.cfg_clk_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05313__B (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05314__A (.DIODE(\u_ws281x.cfg_clk_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05316__A1 (.DIODE(\u_ws281x.cfg_clk_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05320__B1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05326__A (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__05327__A1 (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05327__C1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__05329__B1 (.DIODE(_01123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05329__B2 (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__05330__A1 (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA__05330__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05330__B1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05331__A1 (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05331__A2 (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__05331__A3 (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05331__B1 (.DIODE(\u_glbl_reg.usb_intr_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05332__A1 (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__05332__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05333__A1 (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05333__A2 (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__05333__A3 (.DIODE(_01119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05333__B1 (.DIODE(\u_glbl_reg.i2cm_intr_ss ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05334__A1 (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__05334__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05345__B1 (.DIODE(_01123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05345__B2 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__05346__A1 (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA__05346__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05346__B1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05357__B1 (.DIODE(_01123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05357__B2 (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05358__A1 (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA__05358__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05358__B1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05369__B1 (.DIODE(_01123_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05369__B2 (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__05370__A1 (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA__05370__A2 (.DIODE(_01124_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05370__B1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05371__A_N (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__05371__B (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__05371__C (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05372__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__05372__B (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05373__B (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05373__C (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__05373__D (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05374__B (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__05375__B (.DIODE(_00589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05376__B (.DIODE(_00589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05378__C (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__05378__D (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05379__B (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__05383__B2 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__05384__A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__05385__B (.DIODE(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05387__B (.DIODE(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05388__B (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05389__A2 (.DIODE(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05389__B2 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05390__A2 (.DIODE(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05391__A2 (.DIODE(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05391__B1 (.DIODE(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05392__B1 (.DIODE(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05393__A2 (.DIODE(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05394__A2 (.DIODE(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05395__A2 (.DIODE(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05395__B1 (.DIODE(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05396__A2 (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05396__B1 (.DIODE(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05397__A2 (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05397__B1 (.DIODE(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__A2 (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05398__B1 (.DIODE(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05400__C1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05406__A2 (.DIODE(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__A2 (.DIODE(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05407__B1 (.DIODE(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05408__A2 (.DIODE(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05408__B1 (.DIODE(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__A2 (.DIODE(\u_ws281x.cfg_th0_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05409__B1 (.DIODE(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05410__A1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05410__B1 (.DIODE(\u_ws281x.u_txd_0.led_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05411__A1 (.DIODE(\u_ws281x.u_txd_0.led_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05412__A (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05415__A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__05416__A (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__05417__B (.DIODE(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05418__A_N (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05418__B (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05419__A2 (.DIODE(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05419__B2 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05420__A2 (.DIODE(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05421__A2 (.DIODE(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05421__B1 (.DIODE(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05422__A2 (.DIODE(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05424__B1 (.DIODE(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05425__A2 (.DIODE(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05426__A2 (.DIODE(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05427__A2 (.DIODE(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05427__B1 (.DIODE(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05428__A2 (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05428__B1 (.DIODE(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__A2 (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05429__B1 (.DIODE(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05430__A2 (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05430__B1 (.DIODE(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05431__A2 (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05432__C1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05438__A2 (.DIODE(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05439__A2 (.DIODE(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05439__B1 (.DIODE(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05440__A2 (.DIODE(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05440__B1 (.DIODE(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05441__A2 (.DIODE(\u_ws281x.cfg_th0_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05441__B1 (.DIODE(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05442__A1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05449__D_N (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05451__A (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__A (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__B (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05452__C (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__05453__B (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__A (.DIODE(\u_timer.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05454__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05460__A2 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__05460__C1 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05461__A1 (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05463__B1 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__05464__A (.DIODE(\u_timer.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05464__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__05464__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__A1_N (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05466__B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__05467__A1 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05469__B1 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__05470__A (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__05470__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__05471__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__05473__A1_N (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05473__B1 (.DIODE(net567));
 sky130_fd_sc_hd__diode_2 ANTENNA__05474__A1 (.DIODE(_01332_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A1 (.DIODE(\u_timer.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A2 (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05476__A3 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__05477__B1 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__05479__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05484__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05485__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05486__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05487__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05487__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05488__A1_N (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05488__B2 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05489__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05489__B2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__A1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05490__B2 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05491__A1_N (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05491__B2 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05492__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__05492__B2 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05493__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__A1 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05494__B2 (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05495__A1 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05495__B2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05496__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05497__A1_N (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05497__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05498__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__05499__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05499__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05500__A1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05501__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05501__B2 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05502__A1 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05502__B2 (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05503__B2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05504__A1 (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05504__B2 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05508__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05509__A (.DIODE(_01386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05510__B (.DIODE(_01386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__A_N (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__B (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__C (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__05512__D (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__05513__A (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__B (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA__05514__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__B (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__C (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__05515__D (.DIODE(_01390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05516__A1 (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__05517__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05517__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05518__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05519__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05519__C (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05519__D (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05520__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05521__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05522__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05524__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05525__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05526__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05527__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05529__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05530__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05530__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05531__A1_N (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05531__B2 (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05532__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__05532__B2 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05533__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05533__B2 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05535__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05535__B2 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05536__A1 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05537__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05538__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05539__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05540__A1 (.DIODE(_00882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05541__A1 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05541__B2 (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05542__B2 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05543__A1_N (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05543__B2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__05544__B2 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__A1 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05545__B2 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__A1 (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05546__B2 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05547__A1 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05547__B2 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__05548__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05548__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05551__A2 (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05552__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05556__A1 (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__05558__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__05564__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05566__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05567__B (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05568__A (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05569__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05570__A1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05571__B2 (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05572__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05573__A1_N (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05574__B2 (.DIODE(_00900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05575__A1 (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05576__B2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05577__A1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05577__B2 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05578__A1_N (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05579__B2 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05580__A1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05581__B2 (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05582__B2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05584__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__05585__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05588__A2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05589__B (.DIODE(_01460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05592__A (.DIODE(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05593__A1 (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__05593__B1 (.DIODE(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05594__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05595__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05615__A_N (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05616__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05617__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05627__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__05637__A_N (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05638__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05639__B (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_run ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05639__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05649__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__05659__A_N (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05663__B2 (.DIODE(\u_timer.cfg_pulse_1us[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05664__B2 (.DIODE(\u_timer.cfg_pulse_1us[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05667__B2 (.DIODE(\u_timer.cfg_pulse_1us[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05668__B2 (.DIODE(\u_timer.cfg_pulse_1us[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__A (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__B (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__05673__D (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05674__A (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__05675__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05675__B (.DIODE(_01533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05676__A (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05676__B (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__05676__D (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05677__A (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__05677__B (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05678__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__A (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__B (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05679__C (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05680__A (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__05680__B (.DIODE(_01536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05681__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05681__B (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05682__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__05683__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05683__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05683__C (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__05684__B (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05685__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05685__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05685__C (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__05686__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05687__C (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05688__C (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__05689__A (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05690__C (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__A_N (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__B (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__C (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05691__D (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05692__A (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05693__C (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__05694__A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__05694__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05694__C (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__05695__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05695__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05695__C (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__05696__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05696__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05696__C (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__05697__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05697__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05697__C (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05698__C (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05699__C (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__05700__A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__05700__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05700__C (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__05701__C (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05702__C (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05703__C (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05704__C (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05705__C (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05706__C (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__B (.DIODE(net1177));
 sky130_fd_sc_hd__diode_2 ANTENNA__05707__C (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__B (.DIODE(net1176));
 sky130_fd_sc_hd__diode_2 ANTENNA__05708__C (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05709__C (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__05710__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__05710__B (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA__05710__C (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__B (.DIODE(net1175));
 sky130_fd_sc_hd__diode_2 ANTENNA__05711__C (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__A (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__05712__C (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05713__A (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05713__B (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__A (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05714__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__05715__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05715__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05715__C (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__05716__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05716__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05716__C (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05717__C (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__B (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__05718__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05719__C (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05720__C (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05721__C (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__05722__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05723__C (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__05724__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05724__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05724__C (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__05725__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05725__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05725__C (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__B (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__05726__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05727__C (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05728__C (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05729__C (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__05730__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05730__B (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__05731__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05731__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05731__C (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__05732__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05732__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05732__C (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__05733__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05733__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05733__C (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05734__C (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05735__C (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05736__C (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__05737__A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05737__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05737__C (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05738__C (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05739__C (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__05740__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05740__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05740__C (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__05741__A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05741__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05741__C (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__05742__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05742__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05742__C (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__05743__A (.DIODE(net1319));
 sky130_fd_sc_hd__diode_2 ANTENNA__05743__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05744__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05744__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05744__C (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__05745__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05745__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05745__C (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__05746__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__05746__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05746__C (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__05747__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05747__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05747__C (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__05748__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05748__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05748__C (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__05749__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05749__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05749__C (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__05750__B (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__B (.DIODE(net1173));
 sky130_fd_sc_hd__diode_2 ANTENNA__05751__C (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__05752__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05752__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05752__C (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__05753__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__05753__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05753__C (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__05754__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05754__C (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__05755__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05755__B (.DIODE(net1172));
 sky130_fd_sc_hd__diode_2 ANTENNA__05755__C (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__05756__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05756__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05756__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__05757__A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05757__B (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA__05757__C (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__05758__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05758__C (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__05759__A (.DIODE(net1316));
 sky130_fd_sc_hd__diode_2 ANTENNA__05759__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05759__C (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__A (.DIODE(net1324));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05760__C (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05761__C (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__05762__B (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__05762__C (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05763__C (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__A (.DIODE(net1323));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__B (.DIODE(net1169));
 sky130_fd_sc_hd__diode_2 ANTENNA__05764__C (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__A (.DIODE(net1331));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__B (.DIODE(net1167));
 sky130_fd_sc_hd__diode_2 ANTENNA__05765__C (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__05766__A (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA__05766__B (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__05766__C (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__05767__C (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__05768__C (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__05769__C (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__A_N (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__B_N (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__C (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05770__D (.DIODE(_01003_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05771__C (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__B (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA__05772__C (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05773__C (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05774__C (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05775__C (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05776__C (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__05777__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05777__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05777__C (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05778__C (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__05779__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05779__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05779__C (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05780__C (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__A (.DIODE(net1308));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__B (.DIODE(net1166));
 sky130_fd_sc_hd__diode_2 ANTENNA__05781__C (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05782__C (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__05783__A (.DIODE(net1309));
 sky130_fd_sc_hd__diode_2 ANTENNA__05783__B (.DIODE(net1168));
 sky130_fd_sc_hd__diode_2 ANTENNA__05783__C (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__B (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA__05784__C (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__05785__A (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__05785__B (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05786__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05786__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05786__C (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05787__B (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05788__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__05789__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05789__B (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__05789__C (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05790__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05790__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__05790__C (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05791__A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__05791__B (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA__05791__C (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05792__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05792__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05792__C (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05793__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05793__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__05793__C (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__B (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA__05794__C (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__05795__A (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__05795__B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__05795__C (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__05796__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05796__B (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__05796__C (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__05797__A_N (.DIODE(\u_timer.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05797__C (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__05798__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05798__B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05799__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05799__B (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__05799__C (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__B (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05800__C (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__05801__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05801__B (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA__05801__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__B (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA__05802__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05803__A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA__05803__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__05803__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05804__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05804__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05804__C (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05805__C (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__05806__A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__05806__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__05806__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05807__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__05807__B (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__05807__C (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__B (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__05808__C (.DIODE(net679));
 sky130_fd_sc_hd__diode_2 ANTENNA__05809__A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__05809__B (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__05809__C (.DIODE(net678));
 sky130_fd_sc_hd__diode_2 ANTENNA__05810__A (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__05810__B (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA__05810__C (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__05811__A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__05811__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__05811__C_N (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__05811__D_N (.DIODE(_01002_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05812__A1 (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05813__A1 (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05815__A1 (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05816__A (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__05816__B (.DIODE(_01390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05817__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05817__B (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__05818__B (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__A_N (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__B_N (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__C (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA__05819__D (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__05820__A (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__05821__A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__05822__A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__05823__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05824__A (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05825__A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__05825__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05826__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05826__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05827__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05827__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05828__A (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05829__A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__05829__B (.DIODE(_01566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05830__A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__05830__B (.DIODE(_01566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05831__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05831__B (.DIODE(_01566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05832__A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA__05832__B (.DIODE(_01533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05833__A (.DIODE(net1329));
 sky130_fd_sc_hd__diode_2 ANTENNA__05833__B (.DIODE(_01533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05834__A (.DIODE(net1336));
 sky130_fd_sc_hd__diode_2 ANTENNA__05834__B (.DIODE(_01533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05835__A_N (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05835__C (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA__05835__D (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__05836__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05837__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05837__B (.DIODE(_01565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05838__A (.DIODE(net1313));
 sky130_fd_sc_hd__diode_2 ANTENNA__05838__B (.DIODE(_01566_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05839__A (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__05839__B (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05840__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05840__B (.DIODE(_01567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05841__A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__05841__B (.DIODE(_01567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05842__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__05842__B (.DIODE(_01567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05843__A (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05843__B (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05844__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05844__B (.DIODE(_01568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__A (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__05845__B (.DIODE(_01568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05846__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05846__B (.DIODE(_01568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05847__A (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05847__B (.DIODE(_01534_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05848__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05848__B (.DIODE(_01569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05849__A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__05849__B (.DIODE(_01569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05850__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05850__B (.DIODE(_01569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05851__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05852__A (.DIODE(net1327));
 sky130_fd_sc_hd__diode_2 ANTENNA__05853__A (.DIODE(net1334));
 sky130_fd_sc_hd__diode_2 ANTENNA__05854__B (.DIODE(_01118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05855__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05855__B (.DIODE(_01567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05856__A (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA__05856__B (.DIODE(_01568_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05857__A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA__05857__B (.DIODE(_01569_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05858__A (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__05858__B (.DIODE(_01536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05859__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05859__B (.DIODE(_01570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05860__B (.DIODE(_01570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05861__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__05861__B (.DIODE(_01570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05862__A (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05862__B (.DIODE(_01536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05863__A (.DIODE(net1318));
 sky130_fd_sc_hd__diode_2 ANTENNA__05863__B (.DIODE(_01571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05864__B (.DIODE(_01571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__05865__B (.DIODE(_01571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__A (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05866__B (.DIODE(_01536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05867__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__05867__B (.DIODE(_01572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05868__B (.DIODE(_01572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05869__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__05869__B (.DIODE(_01572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05870__A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA__05870__B (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05871__B (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA__05872__B (.DIODE(_01537_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05873__B (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05873__C (.DIODE(_01388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05874__B (.DIODE(_01570_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05875__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05875__B (.DIODE(_01571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05876__A (.DIODE(net1310));
 sky130_fd_sc_hd__diode_2 ANTENNA__05876__B (.DIODE(_01572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05877__A_N (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__05877__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05878__A_N (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05879__A1 (.DIODE(net1377));
 sky130_fd_sc_hd__diode_2 ANTENNA__05879__A2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05879__B2 (.DIODE(\u_gpio.cfg_gpio_out_data[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05880__A_N (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05881__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05881__A2 (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA__05881__B2 (.DIODE(\u_gpio.cfg_gpio_out_data[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05883__A1 (.DIODE(net1399));
 sky130_fd_sc_hd__diode_2 ANTENNA__05883__A2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05885__A1 (.DIODE(net195));
 sky130_fd_sc_hd__diode_2 ANTENNA__05885__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05886__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05888__A1 (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 ANTENNA__05888__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05890__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05891__A1 (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 ANTENNA__05891__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05892__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05892__B (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__05893__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__05893__C_N (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 ANTENNA__05895__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05897__A1 (.DIODE(_01583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05900__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05901__A1 (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 ANTENNA__05902__A1 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05902__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05905__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05906__A1 (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 ANTENNA__05906__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05907__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05909__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05910__B (.DIODE(\u_gpio.cfg_gpio_dir_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05911__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05911__S (.DIODE(\u_gpio.cfg_gpio_out_type[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05912__A0 (.DIODE(net564));
 sky130_fd_sc_hd__diode_2 ANTENNA__05912__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05914__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05915__A1 (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 ANTENNA__05915__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05916__A1 (.DIODE(_01583_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05916__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05918__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05919__A1 (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 ANTENNA__05919__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05920__A1 (.DIODE(_01584_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05923__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05926__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05928__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05929__A1 (.DIODE(net192));
 sky130_fd_sc_hd__diode_2 ANTENNA__05929__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05931__A1 (.DIODE(net1078));
 sky130_fd_sc_hd__diode_2 ANTENNA__05932__A1 (.DIODE(_01588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05932__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05934__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05936__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__A0 (.DIODE(_01609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__A1 (.DIODE(net191));
 sky130_fd_sc_hd__diode_2 ANTENNA__05937__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__A1 (.DIODE(net193));
 sky130_fd_sc_hd__diode_2 ANTENNA__05938__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05941__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05944__A1 (.DIODE(net1079));
 sky130_fd_sc_hd__diode_2 ANTENNA__05945__A1 (.DIODE(net1414));
 sky130_fd_sc_hd__diode_2 ANTENNA__05945__S (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05946__A2 (.DIODE(_00938_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05947__A2 (.DIODE(_00939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__A1 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__05948__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__A0 (.DIODE(_00936_));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__A1 (.DIODE(net1398));
 sky130_fd_sc_hd__diode_2 ANTENNA__05949__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05950__C (.DIODE(\u_glbl_reg.cfg_multi_func_sel[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05951__B1_N (.DIODE(\u_glbl_reg.cfg_multi_func_sel[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05952__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05953__D (.DIODE(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05954__A (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__05954__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__05955__A_N (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__05955__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05956__A_N (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__05956__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05957__A_N (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__05957__B (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__05958__A1 (.DIODE(net1405));
 sky130_fd_sc_hd__diode_2 ANTENNA__05958__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05959__A1 (.DIODE(net1404));
 sky130_fd_sc_hd__diode_2 ANTENNA__05959__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05960__A1 (.DIODE(net1402));
 sky130_fd_sc_hd__diode_2 ANTENNA__05960__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05961__A1 (.DIODE(net1401));
 sky130_fd_sc_hd__diode_2 ANTENNA__05961__S (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05962__A1 (.DIODE(net1415));
 sky130_fd_sc_hd__diode_2 ANTENNA__05962__S (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__05973__A (.DIODE(\u_glbl_reg.cfg_ref_pll_div[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05976__A1 (.DIODE(\u_glbl_reg.cfg_ref_pll_div[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05977__A (.DIODE(\u_glbl_reg.cfg_ref_pll_div[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A0 (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__A1 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__05988__S (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__05989__A_N (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__05989__B (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__A_N (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__05990__B (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__05991__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05991__B (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__A_N (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA__05992__B (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__05993__A_N (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__05993__B (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__05994__A_N (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__05994__B (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__05995__A_N (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__05995__B (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__05996__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05996__B (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__05997__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05997__B (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__05998__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__05998__B (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__05999__A_N (.DIODE(net1204));
 sky130_fd_sc_hd__diode_2 ANTENNA__05999__B (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__06000__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06000__B (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__06001__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06001__B (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__06002__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06002__B (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__A_N (.DIODE(net1203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06003__B (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__06004__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06004__B (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__06005__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06005__B (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__06006__B (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__06007__B (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__06008__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06008__B (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__06009__B (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06010__B (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__06011__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06011__B (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__06012__A (.DIODE(_00795_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06012__B (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__06013__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06013__A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__06014__A1 (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06014__A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__06015__A1 (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__06015__A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__06016__A1 (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__06016__A2 (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__06017__A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06017__A1 (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__06018__A0 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06018__A1 (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__06027__C (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06029__A (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06042__B1 (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06052__A1 (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__06052__A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__06052__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__A1 (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__06053__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__A1 (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__06054__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06055__A1 (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__06055__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__06055__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06056__A1 (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__06056__A2 (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__06056__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06057__A1 (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__06057__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__06057__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06058__A (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__06058__B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__06059__A1 (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__06059__A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__06059__B1 (.DIODE(\u_glbl_reg.reg_12[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06059__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__A1 (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__B1 (.DIODE(\u_glbl_reg.reg_12[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06060__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06061__A1 (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__06061__A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__06061__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__A1 (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__B1 (.DIODE(\u_glbl_reg.reg_12[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06062__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__A1 (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__B1 (.DIODE(\u_glbl_reg.reg_12[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06063__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__A1 (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__B1 (.DIODE(\u_glbl_reg.reg_12[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06064__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06065__A1 (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__06065__A2 (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__06065__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__A1 (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__A2 (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__B1 (.DIODE(\u_glbl_reg.reg_12[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06066__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06067__A1 (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__06067__B1 (.DIODE(\u_glbl_reg.reg_12[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06067__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__A1 (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__A2 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06068__B1 (.DIODE(\u_glbl_reg.reg_12[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06069__A1 (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__06069__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__A1 (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__A2 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06070__B1 (.DIODE(\u_glbl_reg.reg_12[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06071__A1 (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06071__A2 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06072__A1 (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06072__A2 (.DIODE(_00796_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06072__B1 (.DIODE(\u_glbl_reg.reg_12[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__A1 (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__B1 (.DIODE(\u_glbl_reg.reg_12[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06073__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06074__A (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06075__A1 (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06075__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06075__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__A1 (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__06076__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__A1 (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06077__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06078__A1 (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__06078__A2 (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__06078__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A1 (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__A2 (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06079__B2 (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA__06080__A1 (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__06080__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06080__B2 (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA__06081__A1 (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__06081__B1 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06082__A1 (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA__06082__B1 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06083__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06083__B (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06086__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06086__A2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06086__B1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06087__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06087__B (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06087__C (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06091__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06091__B (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06091__C (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06092__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06093__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06097__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06098__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06101__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06103__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06103__B (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06106__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06106__A2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06106__B1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06110__A (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06113__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06115__A1 (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__06116__S (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06117__A1 (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__06117__S (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06118__A2 (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__06118__S0 (.DIODE(\u_glbl_reg.cfg_mon_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06119__A1 (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA__06119__S0 (.DIODE(\u_glbl_reg.cfg_mon_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06123__A (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__06123__B (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06124__A (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__06125__B (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06126__B (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__A_N (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06127__B (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__06128__B (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__06129__B (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__06130__B (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__A1 (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06131__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06132__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__A2 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06133__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06134__B1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__A2 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06135__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06136__B1 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06137__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06138__B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06140__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06141__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06141__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06142__A2 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06142__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06143__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06143__B1 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06144__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06144__B1 (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA__06145__A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__06145__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06146__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06146__B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06147__A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06147__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06149__A1 (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06149__A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__06149__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06150__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06150__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06151__A2 (.DIODE(_01538_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06151__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06152__B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06153__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06153__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06154__A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06154__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06155__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06156__A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06157__B (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA__06157__C (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06158__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06159__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06159__B1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06160__A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06160__B1 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06162__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06163__A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06163__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06164__A2 (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA__06164__B1 (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06165__A2 (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06166__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06167__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06167__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06168__A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06168__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__06169__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06169__B1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06170__A2 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06170__B1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__06171__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06171__B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06172__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06172__B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06173__A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06173__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06175__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06175__B1 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06176__A2 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06176__B1 (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA__06177__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06177__B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06178__A2 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06178__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06180__A2 (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA__06180__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06181__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06181__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06182__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06183__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06183__B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06184__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06184__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06185__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06185__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06186__A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06186__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__06187__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06187__B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06188__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06188__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06189__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06189__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06190__A2 (.DIODE(net664));
 sky130_fd_sc_hd__diode_2 ANTENNA__06190__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__06191__A2 (.DIODE(net716));
 sky130_fd_sc_hd__diode_2 ANTENNA__06191__B1 (.DIODE(net668));
 sky130_fd_sc_hd__diode_2 ANTENNA__06192__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06192__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__06193__A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06193__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06194__B1 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06195__A2 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06195__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06197__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06197__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06198__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06198__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06199__A2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__06199__B1 (.DIODE(net1137));
 sky130_fd_sc_hd__diode_2 ANTENNA__06200__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06200__B1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06201__A1 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06201__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06201__B1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__06202__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06202__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06202__B2 (.DIODE(\u_gpio.cfg_gpio_dir_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06203__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06203__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06204__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__A1 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06205__B1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__06206__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06206__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06206__B2 (.DIODE(\u_gpio.cfg_gpio_dir_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06207__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06208__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06208__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06209__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06209__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06210__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06211__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06211__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06212__A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__06212__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06213__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06213__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06214__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06214__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06215__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06215__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06216__A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__06216__B1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06217__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06217__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__A1 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06218__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06219__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06219__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06219__B2 (.DIODE(\u_gpio.cfg_gpio_out_data[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06220__A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__06220__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06221__A2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__06221__B1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06222__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06223__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06223__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06223__B2 (.DIODE(\u_gpio.cfg_gpio_out_data[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06224__A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__06224__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06225__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06225__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06226__A2 (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA__06226__B1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06227__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06227__B1 (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__A2 (.DIODE(net717));
 sky130_fd_sc_hd__diode_2 ANTENNA__06228__B1 (.DIODE(net671));
 sky130_fd_sc_hd__diode_2 ANTENNA__06229__A2 (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__06229__B1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__06230__A2 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__06230__B1 (.DIODE(net661));
 sky130_fd_sc_hd__diode_2 ANTENNA__06231__A2 (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__06231__B1 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__06232__A2 (.DIODE(net718));
 sky130_fd_sc_hd__diode_2 ANTENNA__06233__A1 (.DIODE(\u_gpio.u_bit[24].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06233__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06233__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06234__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06235__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06235__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06236__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06237__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06237__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__A1 (.DIODE(net1922));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06238__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06239__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06240__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06240__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06241__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06242__A1 (.DIODE(\u_gpio.u_bit[26].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06242__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06242__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06243__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06243__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06244__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06244__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06245__B1 (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__A1 (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06246__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06247__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06248__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06249__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06249__B1 (.DIODE(net1138));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06250__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06251__B2 (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06252__A2 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06252__B1 (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__A2 (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA__06254__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__A1 (.DIODE(\u_gpio.u_bit[29].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06255__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06256__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06257__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06258__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06258__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06259__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06259__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06260__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06260__B1 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__A2 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06261__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06263__A1 (.DIODE(\u_gpio.cfg_gpio_out_type[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06263__A2 (.DIODE(net702));
 sky130_fd_sc_hd__diode_2 ANTENNA__06263__B1 (.DIODE(net659));
 sky130_fd_sc_hd__diode_2 ANTENNA__06264__A1 (.DIODE(\u_gpio.u_bit[31].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06264__A2 (.DIODE(net691));
 sky130_fd_sc_hd__diode_2 ANTENNA__06264__B1 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06264__B2 (.DIODE(\u_gpio.cfg_gpio_dir_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__A2 (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA__06265__B1 (.DIODE(net1136));
 sky130_fd_sc_hd__diode_2 ANTENNA__06266__A2 (.DIODE(net715));
 sky130_fd_sc_hd__diode_2 ANTENNA__06266__B1 (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__06267__B (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__A1 (.DIODE(\u_glbl_reg.reg_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06268__B2 (.DIODE(\u_glbl_reg.reg_12[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06269__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06269__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__06269__B2 (.DIODE(\u_glbl_reg.cfg_ref_pll_div[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06270__A2 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__06270__B1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__06270__B2 (.DIODE(_01118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__B (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA__06271__C (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__B2 (.DIODE(net2317));
 sky130_fd_sc_hd__diode_2 ANTENNA__06272__C1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__B (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06273__C (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__06274__A (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06274__B (.DIODE(_01118_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__A1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__06277__B2 (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA__06278__A (.DIODE(_01115_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06278__B (.DIODE(_01145_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06279__A1 (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA__06279__A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__06279__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06279__B2 (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 ANTENNA__06279__C1 (.DIODE(_01792_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06280__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06280__B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06281__A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06281__B1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06281__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06282__B (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06283__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06284__A1 (.DIODE(\u_glbl_reg.reg_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06284__B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06285__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06285__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06285__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06288__B (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06289__B (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06290__B (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06294__B2 (.DIODE(\u_glbl_reg.reg_12[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__A2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06295__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__A2 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06296__B2 (.DIODE(net170));
 sky130_fd_sc_hd__diode_2 ANTENNA__06297__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06297__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06298__B1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06299__A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06299__B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06300__A1 (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA__06300__A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06300__B1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06301__B2 (.DIODE(net1099));
 sky130_fd_sc_hd__diode_2 ANTENNA__06302__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06302__A2 (.DIODE(_01805_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06302__A3 (.DIODE(_01807_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06302__B1 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06303__B1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__A1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06304__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06305__A (.DIODE(_01812_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06306__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06306__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06307__A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06307__B1 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06307__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06308__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06308__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06308__B1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06309__B2 (.DIODE(net181));
 sky130_fd_sc_hd__diode_2 ANTENNA__06310__A1 (.DIODE(\u_glbl_reg.reg_2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06310__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06311__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06312__B1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06313__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A1 (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__06320__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__A1 (.DIODE(\u_glbl_reg.reg_23[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__B2 (.DIODE(net1098));
 sky130_fd_sc_hd__diode_2 ANTENNA__06321__C1 (.DIODE(_01833_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06322__B2 (.DIODE(_01832_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06323__A (.DIODE(_01827_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06325__B (.DIODE(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06326__B (.DIODE(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06329__B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06330__A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06330__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06331__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06331__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06331__B2 (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06332__A2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06332__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06332__B2 (.DIODE(\u_glbl_reg.reg_12[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06333__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06333__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06333__B2 (.DIODE(net184));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__A1 (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__06334__B2 (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06335__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06335__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06335__C1 (.DIODE(_01845_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06336__B1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06337__A1 (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA__06337__A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06337__B1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06338__B2 (.DIODE(net1097));
 sky130_fd_sc_hd__diode_2 ANTENNA__06339__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__A2 (.DIODE(_01839_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__A3 (.DIODE(_01840_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06340__B1 (.DIODE(_01851_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06341__A (.DIODE(_01848_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06343__B (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06344__B (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06347__B1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06348__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06349__B2 (.DIODE(net185));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06350__B2 (.DIODE(net1096));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06351__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__A2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06352__B2 (.DIODE(\u_glbl_reg.reg_12[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06353__A1 (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA__06353__A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__06353__B1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__06354__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__06355__A1 (.DIODE(\u_glbl_reg.cfg_mon_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06355__A2 (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA__06355__B1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06356__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06357__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06357__B1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06358__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06358__C1 (.DIODE(_01868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__A1 (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__A2 (.DIODE(_01858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__B1 (.DIODE(_01860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06359__C1 (.DIODE(_01869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06360__B (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06361__B (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06363__B (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06364__B1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06365__A2 (.DIODE(_01857_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06366__B1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__A1 (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__06367__B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06368__B2 (.DIODE(\u_glbl_reg.reg_12[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06369__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06370__B1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__06371__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__A2 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__B2 (.DIODE(net1095));
 sky130_fd_sc_hd__diode_2 ANTENNA__06372__C1 (.DIODE(_01877_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06373__B2 (.DIODE(net186));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06374__B2 (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06375__A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06375__B1 (.DIODE(_01883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06376__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06376__B1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06377__A (.DIODE(_01875_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06378__B (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06379__B (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06381__B (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06382__A2 (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06385__B2 (.DIODE(net1094));
 sky130_fd_sc_hd__diode_2 ANTENNA__06386__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06386__B1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06387__A2 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06388__A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06388__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__A2 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__06389__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06390__B1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06391__B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06392__B2 (.DIODE(net187));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__A1 (.DIODE(net2091));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06393__C1 (.DIODE(_01901_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__A1 (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06394__B1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06395__B1 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06396__C (.DIODE(_01904_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06397__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06397__A2 (.DIODE(_01893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06398__B (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06399__B (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06402__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A1 (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__A2 (.DIODE(net682));
 sky130_fd_sc_hd__diode_2 ANTENNA__06404__B1 (.DIODE(net608));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__A2 (.DIODE(net625));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06405__B2 (.DIODE(\u_glbl_reg.reg_12[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06406__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06407__B1 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__A2 (.DIODE(net655));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06408__B2 (.DIODE(net188));
 sky130_fd_sc_hd__diode_2 ANTENNA__06409__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06410__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06410__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06411__B1 (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06412__B1 (.DIODE(net650));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06413__B2 (.DIODE(net1093));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__A1 (.DIODE(net2097));
 sky130_fd_sc_hd__diode_2 ANTENNA__06414__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__A (.DIODE(_01911_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06415__B (.DIODE(_01919_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06416__B (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__06417__B (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__06419__B (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06420__A2 (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__A (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06422__B (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__A1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__A2 (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06423__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__06424__B2 (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__A2 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06425__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06426__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__A1 (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06427__B1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06428__C1 (.DIODE(_01931_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06429__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06429__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__06430__B2 (.DIODE(net189));
 sky130_fd_sc_hd__diode_2 ANTENNA__06431__A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__06431__B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06432__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06432__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06433__C1 (.DIODE(_01939_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06434__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06435__B1 (.DIODE(_01937_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06436__B (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__06437__B (.DIODE(\u_glbl_reg.u_random.n0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06439__A1 (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06439__A2 (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06441__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06442__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__A2 (.DIODE(net1131));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06443__C1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__A2 (.DIODE(_01550_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06444__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A1 (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06445__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06446__A2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06446__B1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06447__B2 (.DIODE(net190));
 sky130_fd_sc_hd__diode_2 ANTENNA__06448__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06448__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06448__B1 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06449__B2 (.DIODE(\u_glbl_reg.reg_12[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06450__B2 (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06453__A2 (.DIODE(_01946_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06454__B (.DIODE(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06455__B (.DIODE(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06458__A (.DIODE(_01925_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06459__A (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06461__A (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__A2 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06463__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__B1 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06464__C1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06466__A2 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06466__B1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06467__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__A1 (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06468__B2 (.DIODE(\u_glbl_reg.reg_12[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06469__B1 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06470__B2 (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__A1 (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06471__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06472__B1 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06473__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06475__D_N (.DIODE(_01967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06476__B (.DIODE(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06477__B (.DIODE(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06481__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06482__B1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06483__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__A1 (.DIODE(\u_glbl_reg.cfg_rst_ctrl[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06484__B2 (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06485__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A1 (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__A2 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06486__B1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06487__B2 (.DIODE(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06488__B2 (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 ANTENNA__06489__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06490__A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06491__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06492__A2 (.DIODE(_01984_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06493__B (.DIODE(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06494__B (.DIODE(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06500__A1 (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__A2 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06502__B2 (.DIODE(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__A2 (.DIODE(net621));
 sky130_fd_sc_hd__diode_2 ANTENNA__06503__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__A2 (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA__06504__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06505__B1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06506__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06506__B1 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06507__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06508__B2 (.DIODE(net162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__B1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06509__B2 (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__A2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06510__B2 (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06511__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06512__D (.DIODE(_02014_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06513__A2 (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06514__A2 (.DIODE(_02004_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06515__B (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06516__B (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06517__B (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06520__B1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__06522__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A1 (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__A2 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06523__B1 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06524__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06525__B1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06526__B2 (.DIODE(net163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06527__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06528__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06528__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06529__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06530__A2 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06530__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06530__B2 (.DIODE(\u_glbl_reg.reg_12[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__06531__B2 (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA__06532__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06533__A (.DIODE(_02023_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06534__B (.DIODE(net1909));
 sky130_fd_sc_hd__diode_2 ANTENNA__06535__B (.DIODE(\u_glbl_reg.u_random.n0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__A2 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06540__B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__06541__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__A1 (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06542__B1 (.DIODE(net596));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06543__C1 (.DIODE(_02043_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06544__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06545__B1 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06546__B2 (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A1 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__A2 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06547__B2 (.DIODE(net164));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06548__A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06549__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06549__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06550__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A2 (.DIODE(_02039_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__A3 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06551__C1 (.DIODE(_02051_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06555__A2 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__A2 (.DIODE(_02040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06556__B1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__A2 (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA__06558__B1 (.DIODE(net597));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__A2 (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA__06559__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A1 (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__A2 (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06560__B1 (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06561__B1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06562__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__B1 (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA__06563__B2 (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA__06564__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__A2 (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06565__B2 (.DIODE(net165));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__A2 (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06566__B2 (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06567__A2 (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__B1 (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA__06568__C1 (.DIODE(_02067_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06569__A (.DIODE(_02057_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06575__A1 (.DIODE(_01928_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06576__B (.DIODE(net1917));
 sky130_fd_sc_hd__diode_2 ANTENNA__06577__B (.DIODE(\u_glbl_reg.u_random.n0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06579__A (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06580__A (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__06581__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A1 (.DIODE(\u_glbl_reg.reg_2[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__A2 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__B1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06582__C1 (.DIODE(_02080_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06583__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06584__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A1 (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06585__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06586__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06587__B1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__A2 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06588__B2 (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__06589__B2 (.DIODE(net166));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06590__B1 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__A1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06593__B1 (.DIODE(_02091_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06594__B (.DIODE(net1884));
 sky130_fd_sc_hd__diode_2 ANTENNA__06595__B (.DIODE(\u_glbl_reg.u_random.n0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06597__A1 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06599__B2 (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06600__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06601__B1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__B1 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06602__B2 (.DIODE(\u_glbl_reg.reg_2[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__A2 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06603__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__A2 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06604__D1 (.DIODE(_02101_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06605__B1 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__06606__A2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A1 (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06607__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__A2 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06608__C1 (.DIODE(_02105_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06609__D (.DIODE(_02106_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06610__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06611__B (.DIODE(net1931));
 sky130_fd_sc_hd__diode_2 ANTENNA__06612__B (.DIODE(net1931));
 sky130_fd_sc_hd__diode_2 ANTENNA__06616__A (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06619__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__A2 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06620__B2 (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06621__B2 (.DIODE(net168));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06622__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A1 (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06623__B1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__B1 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__06624__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06625__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__A1 (.DIODE(\u_glbl_reg.reg_2[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__A2 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__06626__B1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06627__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06628__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06629__B (.DIODE(_02119_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__A1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06630__B1 (.DIODE(_02126_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06631__B (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__06632__B (.DIODE(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06635__B1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__A2 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__06636__B2 (.DIODE(net169));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06637__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06638__B2 (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06639__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__A1 (.DIODE(\u_glbl_reg.reg_2[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__B1 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06640__B2 (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06641__C1 (.DIODE(_02136_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__A (.DIODE(net1343));
 sky130_fd_sc_hd__diode_2 ANTENNA__06642__C (.DIODE(net1139));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__A2 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06643__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06644__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06644__B1 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__06645__B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__A1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__A2 (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA__06647__B1 (.DIODE(_02133_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06648__B1 (.DIODE(_02143_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06649__B (.DIODE(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06650__B (.DIODE(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06656__A1 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06659__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A1 (.DIODE(\u_glbl_reg.reg_2[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__A2 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__06660__B1 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06661__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06662__A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06663__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A1 (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06664__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__06665__B2 (.DIODE(net171));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__A2 (.DIODE(net700));
 sky130_fd_sc_hd__diode_2 ANTENNA__06666__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06667__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06668__B2 (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA__06669__C (.DIODE(_02161_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06670__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06671__B (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06672__B (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06673__B (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__B1 (.DIODE(net592));
 sky130_fd_sc_hd__diode_2 ANTENNA__06677__B2 (.DIODE(net172));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__A2 (.DIODE(net643));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__B2 (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA__06678__C1 (.DIODE(_02171_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06679__B1 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__06680__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A1 (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06681__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__A1 (.DIODE(\u_glbl_reg.reg_2[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06682__B1 (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA__06683__A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06683__B1 (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA__06684__A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__A2 (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06685__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06686__A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06687__C1 (.DIODE(_02176_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06688__A1 (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA__06689__B (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__06690__B (.DIODE(\u_glbl_reg.u_random.n0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06696__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__A2 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06697__B1 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__A2 (.DIODE(net652));
 sky130_fd_sc_hd__diode_2 ANTENNA__06698__B1 (.DIODE(net614));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B1 (.DIODE(net630));
 sky130_fd_sc_hd__diode_2 ANTENNA__06699__B2 (.DIODE(\u_glbl_reg.reg_22[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A1 (.DIODE(\u_glbl_reg.reg_2[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__A2 (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA__06700__B1 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A1 (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06701__B1 (.DIODE(net610));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A1 (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__A2 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06702__B2 (.DIODE(net173));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__A2 (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA__06703__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06704__A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__A2 (.DIODE(net640));
 sky130_fd_sc_hd__diode_2 ANTENNA__06705__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06706__A2 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06707__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06708__B (.DIODE(\u_glbl_reg.u_random.n0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06709__B (.DIODE(net1905));
 sky130_fd_sc_hd__diode_2 ANTENNA__06712__B1 (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A1 (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__A2 (.DIODE(net684));
 sky130_fd_sc_hd__diode_2 ANTENNA__06713__B1 (.DIODE(net626));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__A2 (.DIODE(net701));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B1 (.DIODE(net562));
 sky130_fd_sc_hd__diode_2 ANTENNA__06714__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__A2 (.DIODE(net639));
 sky130_fd_sc_hd__diode_2 ANTENNA__06715__B1 (.DIODE(net618));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__A2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__B1 (.DIODE(net605));
 sky130_fd_sc_hd__diode_2 ANTENNA__06716__B2 (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__A2 (.DIODE(net1127));
 sky130_fd_sc_hd__diode_2 ANTENNA__06717__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06718__A2 (.DIODE(net635));
 sky130_fd_sc_hd__diode_2 ANTENNA__06719__A2 (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__A2 (.DIODE(net623));
 sky130_fd_sc_hd__diode_2 ANTENNA__06720__B1 (.DIODE(net611));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A1 (.DIODE(\u_glbl_reg.reg_15[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__A2 (.DIODE(net657));
 sky130_fd_sc_hd__diode_2 ANTENNA__06721__B1 (.DIODE(net647));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A1 (.DIODE(\u_glbl_reg.reg_2[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__A2 (.DIODE(net687));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__B1 (.DIODE(net591));
 sky130_fd_sc_hd__diode_2 ANTENNA__06722__B2 (.DIODE(net174));
 sky130_fd_sc_hd__diode_2 ANTENNA__06723__C (.DIODE(_02214_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06725__B (.DIODE(\u_glbl_reg.u_random.n0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06726__B (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__06732__A1 (.DIODE(_02074_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06734__B1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A1 (.DIODE(\u_glbl_reg.reg_2[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06735__B1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06736__B1 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06737__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06738__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A1 (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06739__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__A2 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06740__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06741__B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06742__B2 (.DIODE(net1107));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06743__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06745__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06746__B1 (.DIODE(_02236_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06747__B (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06748__B (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06752__A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__A1 (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06753__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__A1 (.DIODE(\u_glbl_reg.reg_2[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__B1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06754__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06755__B1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06756__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06757__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06758__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06759__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__B2 (.DIODE(net1106));
 sky130_fd_sc_hd__diode_2 ANTENNA__06760__C1 (.DIODE(_02249_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06761__B1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06762__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06763__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06764__A (.DIODE(_02242_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06765__B (.DIODE(net1915));
 sky130_fd_sc_hd__diode_2 ANTENNA__06766__B (.DIODE(net1915));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__A2 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__06771__B1 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06772__B1 (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06773__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06774__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06775__B2 (.DIODE(net1105));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__B1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06776__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06777__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06778__B1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06779__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06780__A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06781__B (.DIODE(_02265_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06782__C (.DIODE(_02270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06783__B1 (.DIODE(_02271_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06784__B (.DIODE(net1894));
 sky130_fd_sc_hd__diode_2 ANTENNA__06785__B (.DIODE(net1894));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06788__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06789__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__B1 (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA__06790__B2 (.DIODE(net1104));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06791__B1 (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA__06792__A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A1 (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06793__B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A1 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06794__B2 (.DIODE(net178));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06795__B1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06796__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06797__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__A1 (.DIODE(net593));
 sky130_fd_sc_hd__diode_2 ANTENNA__06799__B1 (.DIODE(_02286_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06807__A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06808__B1 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06809__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06810__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06811__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06812__A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A1 (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06813__B1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__A2 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__B1 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06814__B2 (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A1 (.DIODE(\u_glbl_reg.reg_2[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06815__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06816__B2 (.DIODE(net1103));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06817__B2 (.DIODE(net179));
 sky130_fd_sc_hd__diode_2 ANTENNA__06819__B1 (.DIODE(_02305_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06820__B (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06821__B (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__A2 (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA__06825__B1 (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__A2 (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06826__B2 (.DIODE(net1102));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__A2 (.DIODE(net698));
 sky130_fd_sc_hd__diode_2 ANTENNA__06827__B1 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06828__B1 (.DIODE(net645));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06829__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__A1 (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06830__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06831__B1 (.DIODE(net589));
 sky130_fd_sc_hd__diode_2 ANTENNA__06832__A2 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06833__B1 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__B1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__B2 (.DIODE(_02310_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06834__C1 (.DIODE(_02319_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06835__A2 (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA__06836__B (.DIODE(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06837__B (.DIODE(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06839__B2 (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06842__A (.DIODE(_01789_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__A2 (.DIODE(net624));
 sky130_fd_sc_hd__diode_2 ANTENNA__06843__B1 (.DIODE(net612));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__A2 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06844__B1 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A1 (.DIODE(\u_glbl_reg.reg_2[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06845__B1 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06846__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06847__B1 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__A2 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06848__B1 (.DIODE(net607));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__A2 (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__B1 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06849__B2 (.DIODE(net1101));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__B1 (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA__06850__B2 (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06851__B2 (.DIODE(net182));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__A2 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06852__B2 (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__06854__A (.DIODE(_02327_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06856__B (.DIODE(\u_glbl_reg.u_random.n0[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__A2 (.DIODE(net620));
 sky130_fd_sc_hd__diode_2 ANTENNA__06858__B1 (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__A2 (.DIODE(net641));
 sky130_fd_sc_hd__diode_2 ANTENNA__06859__B1 (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__A2 (.DIODE(net1124));
 sky130_fd_sc_hd__diode_2 ANTENNA__06860__B1 (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__A1 (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__A2 (.DIODE(net681));
 sky130_fd_sc_hd__diode_2 ANTENNA__06861__B1 (.DIODE(net628));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__A1 (.DIODE(\u_glbl_reg.reg_2[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__A2 (.DIODE(net685));
 sky130_fd_sc_hd__diode_2 ANTENNA__06862__B1 (.DIODE(net654));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A1 (.DIODE(net1100));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__A2 (.DIODE(net603));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B1 (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA__06863__B2 (.DIODE(net183));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__A2 (.DIODE(net649));
 sky130_fd_sc_hd__diode_2 ANTENNA__06864__B1 (.DIODE(net646));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__A2 (.DIODE(net699));
 sky130_fd_sc_hd__diode_2 ANTENNA__06865__B1 (.DIODE(_01786_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06866__A2 (.DIODE(net637));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__A2 (.DIODE(net633));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__B1 (.DIODE(net616));
 sky130_fd_sc_hd__diode_2 ANTENNA__06867__B2 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06868__A2 (.DIODE(net560));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A1 (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA__06869__A2 (.DIODE(_02341_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06870__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06871__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06872__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06873__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06874__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06875__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06876__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__A1 (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA__06877__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06878__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06879__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06880__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06881__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06882__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06883__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06884__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06885__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06886__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06887__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__06888__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06889__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06890__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06891__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06892__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06893__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06894__B (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06895__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06896__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06897__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06898__C1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__06899__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06900__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06901__C1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__06902__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06903__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06904__C1 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__06905__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06906__B (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06907__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06908__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06909__B (.DIODE(net1367));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06910__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06911__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06912__B (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__A1 (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06913__C1 (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__06914__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__06915__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06916__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06917__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06918__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06919__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06920__A2 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06921__B (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06922__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06923__A2 (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06924__B (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__B2 (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_2[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06925__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06926__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA__06927__B (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__A1 (.DIODE(net1278));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06928__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06929__A2 (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06930__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__A1 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06931__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06932__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__06933__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__A1 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B1 (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06934__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06935__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06936__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__A1 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06937__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06938__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__A (.DIODE(net1360));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__B (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA__06939__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__A1 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B1 (.DIODE(net1162));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__B2 (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06940__C1 (.DIODE(net1245));
 sky130_fd_sc_hd__diode_2 ANTENNA__06941__A2 (.DIODE(net1229));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06942__B (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__B1 (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA__06943__C1 (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06944__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__A (.DIODE(_00941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06945__B (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__B1 (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA__06946__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06947__B2 (.DIODE(_02404_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06948__B (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06949__C1 (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06950__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06951__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__B1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__06952__C1 (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06953__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06954__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__B1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__06955__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__06956__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06957__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__B1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__06958__C1 (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__06959__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__06960__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06961__C1 (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06962__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__B (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__06963__C (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__B1 (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA__06964__C1 (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA__06965__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06968__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06981__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06982__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06985__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06987__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06989__B (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06990__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06991__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06992__B (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06993__A2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06994__A2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06995__B (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06996__B (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06997__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__06999__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07000__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07002__A2 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07003__A3 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07004__C1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07005__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07006__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07007__B2 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07008__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07009__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A1 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07010__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07011__A1 (.DIODE(_00900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07012__B2 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07013__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07014__A (.DIODE(_00900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__A (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07015__B (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07016__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07017__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07019__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__A (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07020__B (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A1 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07021__B2 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07029__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07032__B2 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07036__A1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07037__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07038__B2 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07040__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07041__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A1 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07043__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__A1 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07044__B2 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__A1_N (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07049__B2 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__07050__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07051__A (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__07053__B1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07054__A (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__A2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07059__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07060__B (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07071__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07073__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07074__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07075__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07077__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07080__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07081__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07082__A2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07085__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07086__B1 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07104__B (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07105__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07106__C (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07110__C1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07111__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07112__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07114__B2 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07120__A1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07122__B2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__A1 (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07123__B2 (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07124__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07125__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__07126__A1 (.DIODE(_00900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07128__A (.DIODE(_00900_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07135__B (.DIODE(_02585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07146__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07147__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07149__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07150__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07151__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07154__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__A2 (.DIODE(_02446_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07155__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07156__B (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__A2 (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07157__B1 (.DIODE(_02447_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07159__C (.DIODE(_02443_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07160__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__07161__B2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07162__B1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07163__B2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__A2_N (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07168__B1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07171__B2 (.DIODE(_00899_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07172__C1 (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07173__A1 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__A1 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07174__B2 (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07175__B2 (.DIODE(_00910_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07176__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07177__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A1 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07178__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__A1 (.DIODE(_00905_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07180__B2 (.DIODE(_00906_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07181__A (.DIODE(_00898_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07182__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07194__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07195__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07196__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07197__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07198__C1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07199__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07200__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07201__C1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07202__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__07203__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07204__C1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07205__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07206__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07207__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07208__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07209__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07210__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07211__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07212__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07213__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07214__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07215__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07216__C1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07217__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07218__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__A2 (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07219__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07220__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07221__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__A2 (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07222__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07223__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07224__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07225__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07226__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07227__C (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07228__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07229__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07230__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07231__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07232__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07233__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07234__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07235__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07236__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07237__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07238__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07239__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07240__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07241__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07242__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07243__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07244__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07245__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07246__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07247__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07248__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07249__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07250__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07251__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07252__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07253__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07254__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__A1 (.DIODE(net1268));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07255__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07256__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__A (.DIODE(net1350));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07257__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07258__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07259__A2 (.DIODE(net1219));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07260__C (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07261__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07262__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07263__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__B2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07264__C1 (.DIODE(net1236));
 sky130_fd_sc_hd__diode_2 ANTENNA__07265__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07266__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07267__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07268__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07269__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07270__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07271__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07272__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07273__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07274__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07275__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07276__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07277__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07278__B (.DIODE(net1362));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07279__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07280__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07281__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07282__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07283__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07284__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__B1 (.DIODE(net1154));
 sky130_fd_sc_hd__diode_2 ANTENNA__07285__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07286__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__A (.DIODE(net1348));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07287__C (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__A1 (.DIODE(net1266));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__B1 (.DIODE(net1142));
 sky130_fd_sc_hd__diode_2 ANTENNA__07288__C1 (.DIODE(net1234));
 sky130_fd_sc_hd__diode_2 ANTENNA__07289__A2 (.DIODE(net1217));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07290__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07291__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07292__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07293__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07294__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07295__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07296__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07297__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07298__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07299__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07300__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07301__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07302__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07303__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07304__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07305__B (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07306__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07307__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07308__B (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07309__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07310__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07311__B (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07312__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07313__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__A (.DIODE(_00961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07314__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07315__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07316__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07317__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07318__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07319__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07320__B (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07321__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07322__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07323__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07324__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07325__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07326__B (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07327__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07328__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07329__B (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07330__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07331__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07332__B (.DIODE(net1212));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07333__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07334__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07335__B (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__A1 (.DIODE(net1273));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07336__C1 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07337__A2 (.DIODE(net1223));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07338__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07339__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07340__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07341__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07342__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07343__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__07344__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07345__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07346__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07347__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07348__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07349__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__07350__B (.DIODE(net1256));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__A1 (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07351__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07352__A2 (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07353__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__A1 (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__B1 (.DIODE(net1155));
 sky130_fd_sc_hd__diode_2 ANTENNA__07354__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07355__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__B (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA__07356__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07357__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07358__A2 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA__07359__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__A1 (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07360__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07361__A2 (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07362__B (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07363__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07364__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07365__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__B1 (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA__07366__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07367__A2 (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__B (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA__07368__C (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__B2 (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__07369__C1 (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA__07370__A2 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__A (.DIODE(_00967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07371__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__A1 (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__B2 (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA__07372__C1 (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA__07373__A2 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__A (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07374__B (.DIODE(net1211));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__B1 (.DIODE(net1156));
 sky130_fd_sc_hd__diode_2 ANTENNA__07375__C1 (.DIODE(net1237));
 sky130_fd_sc_hd__diode_2 ANTENNA__07376__A2 (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__A (.DIODE(_00969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07377__B (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__B2 (.DIODE(net2105));
 sky130_fd_sc_hd__diode_2 ANTENNA__07378__C1 (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA__07379__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07380__B (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07381__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07382__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__A (.DIODE(net1352));
 sky130_fd_sc_hd__diode_2 ANTENNA__07383__B (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B1 (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07384__C1 (.DIODE(net1241));
 sky130_fd_sc_hd__diode_2 ANTENNA__07385__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__07386__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07387__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07388__B (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07392__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07394__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07400__B1 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07403__A2 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07404__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B1 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07405__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07407__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07408__B1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07409__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07410__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07411__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07412__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07413__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07414__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07415__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07417__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__A (.DIODE(net1076));
 sky130_fd_sc_hd__diode_2 ANTENNA__07418__B (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__A2 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07419__B1 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07420__B (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07421__B1 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07425__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07426__A (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07427__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__A1 (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07429__B2 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A1 (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07430__B2 (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A1 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07431__B2 (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07432__B2 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__A1 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07433__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07437__C1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07438__B2 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__A1 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07439__B2 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__A1 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07440__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07441__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__A1 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07442__B2 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07444__B2 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A1 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07445__B2 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07446__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07448__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07451__A1 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__A1 (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07454__B2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07455__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07457__A (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07458__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__A1 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07459__B2 (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07461__B2 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07462__C1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__A1 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07463__B2 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__A1 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07464__B2 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__A1 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07466__B2 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07467__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07469__B2 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__A1 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07470__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A1 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07472__B2 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A1 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07474__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__A1 (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07475__B2 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07477__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__A2 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07478__B1 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07479__B1 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07480__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07481__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07483__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07489__B1 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07491__A2 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07492__B (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07494__B1 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__A2_N (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07495__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07498__A2 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07499__A2 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07500__B2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07503__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07505__A1_N (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07506__A (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07507__C1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__A1 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07508__B2 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__A1 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07509__B2 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__A1 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07511__B2 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07512__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__A1 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07514__B2 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07515__A1 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__A1 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07516__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07518__B (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__A2_N (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07519__B1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07521__B2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__A1 (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07522__B2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07523__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07524__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__A1 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07525__B2 (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07526__A (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07527__A (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07528__A (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__A2 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07532__B1 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07533__B1 (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07534__B1 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07536__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07542__B1 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07544__A2 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07545__B1 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__A2 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07548__B1 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07551__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07552__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07553__B1 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07555__A3 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07560__B (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07561__A (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__A1 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07562__B2 (.DIODE(_00859_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__A1 (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07563__B2 (.DIODE(_00860_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A1_N (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07564__A2_N (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07565__A (.DIODE(_00861_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__A (.DIODE(_00862_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07566__B (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__A1_N (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B1 (.DIODE(_00941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07568__B2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07569__A2 (.DIODE(_00941_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07573__C1 (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__A1 (.DIODE(_00872_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07574__B2 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__A1 (.DIODE(_00871_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07575__B2 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A1 (.DIODE(_00870_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07576__B2 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A1 (.DIODE(_00869_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07577__B2 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A1 (.DIODE(_00868_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07578__B2 (.DIODE(net728));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07579__B2 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07580__B2 (.DIODE(_00863_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A1 (.DIODE(_00866_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__A2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07581__B2 (.DIODE(_00865_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__A (.DIODE(_00858_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07582__B (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07588__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07589__B (.DIODE(_02803_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B1 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07590__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07591__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07592__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07595__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07596__C1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07598__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07600__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B1 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07601__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__A2 (.DIODE(_02785_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07602__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B1 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07603__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__A2 (.DIODE(_02773_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B1 (.DIODE(_02790_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07604__B2 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07605__A2 (.DIODE(_02793_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07607__A2 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07608__B (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__A2 (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07609__B1 (.DIODE(_02804_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07610__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__B (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07611__C (.DIODE(_02799_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07619__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07621__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07622__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07625__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07626__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__A2 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07627__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07629__B1 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07630__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__A2 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07631__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07632__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07635__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07636__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07637__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B1 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07638__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07639__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07641__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07642__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07643__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07644__B (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07645__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07646__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07647__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07648__B (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07649__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07651__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07653__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07654__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07655__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__A (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__07656__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07657__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07658__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07660__B1 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07668__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07670__B2 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07671__B2 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07672__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07673__A (.DIODE(_00882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__A (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07674__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07676__A (.DIODE(_00882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07677__A (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A1 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07678__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__A1 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07681__B2 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__A1 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07682__B2 (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07683__A (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__A (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07684__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07687__B2 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07688__A (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07689__A_N (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07690__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A1_N (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__A2_N (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07693__B1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__A (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07694__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07696__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__A (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07699__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__A (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07700__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__A (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07701__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07702__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07703__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07705__C_N (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07709__A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07712__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07716__A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__A1 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07717__B2 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__A1 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07718__B2 (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07719__A (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__A1 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07720__B2 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07721__A_N (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07722__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07723__A1 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07724__B2 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07725__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07728__A (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07729__A (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__A1 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07731__B2 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07732__A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07733__B2 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07734__A_N (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07735__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07736__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07737__B1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A1 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07738__B2 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__A (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07739__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07740__A1 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07743__A (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07745__A1 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07748__A (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07751__B2 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07756__B (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__A2 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07757__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07758__B1 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__A2 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07759__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07761__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07762__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07763__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07764__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07765__B1 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07766__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07767__B (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07768__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07770__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07771__A2 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07773__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07774__A2 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07778__B (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07779__A2 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07781__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__B1 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07788__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__A2 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07789__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__A2 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07790__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07793__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07795__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07797__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07798__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07799__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07800__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07801__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07802__B (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07803__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B1 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07804__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07815__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07817__A (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A1 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07818__B2 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__A1 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07819__B2 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07821__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__A1_N (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07822__B1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07823__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__A1 (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07824__B2 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__A1 (.DIODE(_00881_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07825__B2 (.DIODE(_00880_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07827__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07829__B2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__A1 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07830__B2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__A1 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07831__B2 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07832__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__A (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07833__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07834__B2 (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07837__B2 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07839__B2 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07842__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__A (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07843__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07845__A2 (.DIODE(_00961_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07848__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07849__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B1 (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07855__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07856__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__A2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B1 (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07857__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07858__B (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B1 (.DIODE(_03022_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07859__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07861__B2 (.DIODE(net588));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07862__B (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07863__B (.DIODE(net587));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07864__A2 (.DIODE(_03030_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__B1 (.DIODE(_03031_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07865__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__A2 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07868__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07870__B1 (.DIODE(_03015_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07871__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B1 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07873__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07874__A2 (.DIODE(_03006_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__A2 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07875__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07878__B (.DIODE(_03027_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__A2 (.DIODE(_03010_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__B1 (.DIODE(_03011_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07880__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07884__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07885__A2 (.DIODE(_03021_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__A (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07888__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A1 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07889__B2 (.DIODE(_00882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A1 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07890__B2 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A1 (.DIODE(_00884_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07891__B2 (.DIODE(_00883_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__A2 (.DIODE(_00969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07893__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__A2 (.DIODE(_00967_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07894__B1 (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A1_N (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__A2_N (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07895__B1 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__A2 (.DIODE(_00968_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B1 (.DIODE(_00969_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07896__B2 (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A1 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07898__B2 (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A1 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07899__B2 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A1 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07900__B2 (.DIODE(_00889_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__A (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07901__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07902__B2 (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07903__B2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A1 (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07904__B2 (.DIODE(_00890_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A1 (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07906__B2 (.DIODE(_00887_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__A (.DIODE(_00886_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07909__B (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A1 (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07910__B2 (.DIODE(net727));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A1 (.DIODE(_00892_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07915__A2 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07916__A1 (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07925__B (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A1 (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__A2 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__07926__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07927__B (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A1 (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__A2 (.DIODE(net1244));
 sky130_fd_sc_hd__diode_2 ANTENNA__07928__B1 (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__A (.DIODE(net1355));
 sky130_fd_sc_hd__diode_2 ANTENNA__07929__B (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__A2 (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07930__B1 (.DIODE(net1157));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__07931__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__A (.DIODE(net1354));
 sky130_fd_sc_hd__diode_2 ANTENNA__07932__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA__07933__B (.DIODE(net1261));
 sky130_fd_sc_hd__diode_2 ANTENNA__07934__B (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__07935__B (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__A (.DIODE(net1826));
 sky130_fd_sc_hd__diode_2 ANTENNA__07936__B (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07937__B (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__07938__B (.DIODE(net1239));
 sky130_fd_sc_hd__diode_2 ANTENNA__07939__B (.DIODE(net1243));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07940__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA__07941__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07942__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA__07943__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07944__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07945__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07946__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07947__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07948__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07949__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07950__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07951__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07952__C1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07953__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07954__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07955__C1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07956__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07957__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA__07958__B (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__07959__C1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__07960__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07961__B (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__07962__C1 (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__07963__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07964__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07965__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A1 (.DIODE(\u_timer.cfg_pulse_1us[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07966__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07967__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07968__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A1 (.DIODE(\u_timer.cfg_pulse_1us[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__07969__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07970__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07971__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07972__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__B1 (.DIODE(net1148));
 sky130_fd_sc_hd__diode_2 ANTENNA__07973__C1 (.DIODE(net1250));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07974__B (.DIODE(net1370));
 sky130_fd_sc_hd__diode_2 ANTENNA__07975__A2 (.DIODE(net1231));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__A (.DIODE(net1282));
 sky130_fd_sc_hd__diode_2 ANTENNA__07976__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07977__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07978__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__07979__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07980__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07981__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__07982__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07983__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07984__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07985__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__07986__B (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__07987__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07988__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__A1 (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07989__B1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__07990__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07991__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__07992__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07993__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__A (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__07994__B (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__A1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__B2 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__07995__C1 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__07996__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07997__B1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__07998__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__07999__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08000__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08001__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08002__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08003__B1 (.DIODE(net1262));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__A1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08004__B1 (.DIODE(net1150));
 sky130_fd_sc_hd__diode_2 ANTENNA__08005__A2 (.DIODE(net1232));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08006__B1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08007__A1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08008__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08009__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08010__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08011__A2 (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__08012__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__08013__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08014__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__08015__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__A1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08016__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08017__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08018__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08019__B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08020__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08021__B1 (.DIODE(net1260));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08022__B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08023__A2 (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08024__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__A1 (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA__08025__B1 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__08026__A2 (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA__08027__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__08028__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08029__A2 (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA__08030__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__A1 (.DIODE(net1271));
 sky130_fd_sc_hd__diode_2 ANTENNA__08031__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08032__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__08033__B1 (.DIODE(net1258));
 sky130_fd_sc_hd__diode_2 ANTENNA__08034__B1 (.DIODE(net1143));
 sky130_fd_sc_hd__diode_2 ANTENNA__08035__A2 (.DIODE(net1222));
 sky130_fd_sc_hd__diode_2 ANTENNA__08036__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08037__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__A2 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08038__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__A1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B1 (.DIODE(_03377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08039__B2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A1 (.DIODE(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08040__B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__08042__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08043__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B1 (.DIODE(_03382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08044__B2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A1 (.DIODE(\u_ws281x.cfg_reset_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08045__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A1 (.DIODE(\u_ws281x.cfg_clk_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__A2 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B1 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08046__B2 (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A1 (.DIODE(\u_ws281x.cfg_clk_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__A2 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__08048__B1 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08049__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08050__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B1 (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08051__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A1 (.DIODE(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08052__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A1 (.DIODE(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08053__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08054__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08055__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__A1 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__08056__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08057__A2 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A1 (.DIODE(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08058__B1 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08059__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08060__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08061__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A1 (.DIODE(\u_ws281x.cfg_clk_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08062__A2 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A1 (.DIODE(\u_ws281x.cfg_clk_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__A2 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B1 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__08063__B2 (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08064__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08065__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08066__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08067__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08068__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08069__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__A2 (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08070__B2 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A1 (.DIODE(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08071__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08072__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08073__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__A2 (.DIODE(_03405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08074__B2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08075__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08076__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08077__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__A2 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08078__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08079__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08080__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08081__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08082__B2 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A1 (.DIODE(\u_ws281x.cfg_reset_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08083__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08084__S (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA__08085__S (.DIODE(net1084));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__A1 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08086__B2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A1 (.DIODE(\u_ws281x.cfg_reset_period[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08087__B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__08088__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08089__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08090__B2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08091__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08092__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08093__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__A1 (.DIODE(net712));
 sky130_fd_sc_hd__diode_2 ANTENNA__08094__B2 (.DIODE(net708));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__A2 (.DIODE(net705));
 sky130_fd_sc_hd__diode_2 ANTENNA__08095__B1 (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA__08096__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08097__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08098__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08099__B1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08100__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08101__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08102__B2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A1 (.DIODE(\u_ws281x.cfg_reset_period[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08103__B1 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08104__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08105__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08106__B2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A1 (.DIODE(\u_ws281x.cfg_reset_period[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__A2 (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA__08107__B1 (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA__08108__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08109__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08110__A2 (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A1 (.DIODE(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08111__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08112__S (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA__08113__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08114__A2 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A1 (.DIODE(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08115__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08116__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__A (.DIODE(_00996_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08117__B (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA__08118__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A1 (.DIODE(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B1 (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08119__B2 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08120__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08121__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08122__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A1 (.DIODE(\u_ws281x.cfg_th0_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08123__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08124__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08125__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__A (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08126__C (.DIODE(_03445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A1 (.DIODE(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08127__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08128__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08129__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08130__B1 (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A1 (.DIODE(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08131__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08132__S (.DIODE(net1080));
 sky130_fd_sc_hd__diode_2 ANTENNA__08133__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__A (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08134__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A1 (.DIODE(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08135__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08136__S (.DIODE(net1083));
 sky130_fd_sc_hd__diode_2 ANTENNA__08137__S (.DIODE(net1081));
 sky130_fd_sc_hd__diode_2 ANTENNA__08138__A1 (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA__08139__A2 (.DIODE(net694));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__A (.DIODE(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08140__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__A (.DIODE(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08141__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__A (.DIODE(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08142__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__A (.DIODE(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08143__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__A (.DIODE(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08144__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__A (.DIODE(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08145__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08146__C (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__B (.DIODE(net1164));
 sky130_fd_sc_hd__diode_2 ANTENNA__08147__C (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA__08148__C_N (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08150__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08151__B2 (.DIODE(_03458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08152__B (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08153__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08154__C (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__B1 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08155__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08156__A_N (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__08157__A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__08158__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08159__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__A2 (.DIODE(\u_timer.reg_rdata[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__B1 (.DIODE(_03463_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08160__C1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08161__B (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__08162__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08163__A (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08164__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__A2 (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA__08165__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08166__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08167__A (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__B (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08170__C (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__A1 (.DIODE(_03473_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08171__B1 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08172__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08173__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08174__B2 (.DIODE(_03480_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08175__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__A2 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08176__C1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__A2 (.DIODE(\u_timer.reg_rdata[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08177__C1 (.DIODE(_03483_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__A2 (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA__08178__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08179__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08180__B1 (.DIODE(_03485_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08181__B2 (.DIODE(_03487_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08182__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08183__B2 (.DIODE(_03488_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08184__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__A2 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08185__C1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08186__C1 (.DIODE(_03491_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__A2 (.DIODE(net88));
 sky130_fd_sc_hd__diode_2 ANTENNA__08187__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08188__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08189__B1 (.DIODE(_03493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08190__B2 (.DIODE(_03495_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08191__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08192__B2 (.DIODE(_03496_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08193__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__A2 (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08194__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08195__C1 (.DIODE(_03499_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__A2 (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA__08196__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08197__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08198__B1 (.DIODE(_03501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08200__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08201__B2 (.DIODE(_03504_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08202__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08203__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08204__C1 (.DIODE(_03507_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08205__A2 (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 ANTENNA__08206__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08207__B1 (.DIODE(_03509_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08208__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08209__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08210__B2 (.DIODE(_03512_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08211__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08212__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08213__C1 (.DIODE(_03515_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08214__A2 (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 ANTENNA__08215__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08216__B1 (.DIODE(_03517_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08217__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__A2 (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 ANTENNA__08218__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08219__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08220__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08221__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08224__C1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__A2 (.DIODE(_03523_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08225__B1 (.DIODE(_03526_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08226__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08227__B1 (.DIODE(_03527_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08228__A2 (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08230__S (.DIODE(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08231__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08232__C1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08233__B1 (.DIODE(_03533_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08234__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08235__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08236__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08237__B2 (.DIODE(_03536_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08238__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08239__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__A2 (.DIODE(\u_timer.reg_rdata[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08240__C1 (.DIODE(_03539_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08241__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08242__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08243__B1 (.DIODE(_03541_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08244__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08245__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__A2 (.DIODE(net1121));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B1 (.DIODE(net1116));
 sky130_fd_sc_hd__diode_2 ANTENNA__08246__B2 (.DIODE(_03544_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08247__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08248__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__A2 (.DIODE(\u_timer.reg_rdata[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08249__C1 (.DIODE(_03547_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08250__A2 (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 ANTENNA__08251__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08252__B1 (.DIODE(_03549_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08253__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08254__B (.DIODE(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08255__B2 (.DIODE(_03552_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08256__B (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08257__C1 (.DIODE(net1092));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A1 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__A2 (.DIODE(\u_timer.reg_rdata[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__B1 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08258__C1 (.DIODE(_03555_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__A2 (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA__08259__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08260__B (.DIODE(net549));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08261__B1 (.DIODE(_03557_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08262__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08263__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08265__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08266__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__B1 (.DIODE(_03560_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08267__C1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08268__B1 (.DIODE(_03564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08269__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08270__B1 (.DIODE(_03565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08271__A2 (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A0 (.DIODE(\u_pwm.reg_rdata_pwm0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08273__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08274__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__B1 (.DIODE(_03567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08275__C1 (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08276__B1 (.DIODE(_03571_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08277__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08278__B1 (.DIODE(_03572_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08279__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__A0 (.DIODE(\u_pwm.reg_rdata_pwm0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08281__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08282__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__B1 (.DIODE(_03574_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08283__C1 (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08284__B1 (.DIODE(_03578_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08285__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08286__B1 (.DIODE(_03579_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08287__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08289__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A1 (.DIODE(\u_pwm.reg_rdata_pwm1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08290__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__B1 (.DIODE(_03581_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08291__C1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08292__B1 (.DIODE(_03585_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08293__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08294__B1 (.DIODE(_03586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08295__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__A1 (.DIODE(\u_pwm.reg_rdata_pwm2[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08297__S (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08298__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__A2 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__B1 (.DIODE(_03588_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08299__C1 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__A2 (.DIODE(_03591_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08300__B1 (.DIODE(_03592_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08301__B (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__A2 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08302__B1 (.DIODE(_03593_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08303__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08304__B2 (.DIODE(_03595_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08305__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08306__B1 (.DIODE(_03596_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__A2 (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA__08307__C1 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__A1 (.DIODE(\u_timer.reg_rdata[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__B1 (.DIODE(_03598_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__B2 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08308__C1 (.DIODE(_03599_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08309__S (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08310__B1 (.DIODE(_03601_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08311__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08312__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08313__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__B1 (.DIODE(_03603_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08314__C1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__A2 (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08315__C1 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__A1 (.DIODE(\u_timer.reg_rdata[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__B1 (.DIODE(_03605_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08316__C1 (.DIODE(_03606_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08317__S (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08318__B1 (.DIODE(_03608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08319__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08320__B2 (.DIODE(_03609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08321__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__B1 (.DIODE(_03610_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08322__C1 (.DIODE(_03467_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__A2 (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA__08323__C1 (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__B1 (.DIODE(_03612_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08324__C1 (.DIODE(_03613_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08325__S (.DIODE(_03476_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08326__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__A2 (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA__08327__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08328__B (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__A2 (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA__08329__B1 (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA__08330__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08331__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08332__A2 (.DIODE(_03618_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__A1 (.DIODE(\u_glbl_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08333__B1 (.DIODE(net1795));
 sky130_fd_sc_hd__diode_2 ANTENNA__08334__A2 (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA__08335__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08336__B2 (.DIODE(_03623_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08337__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08338__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08339__A2 (.DIODE(_03624_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08340__B1 (.DIODE(_03622_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08341__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08342__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08343__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08344__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__A2 (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08345__B1 (.DIODE(net540));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08346__A2 (.DIODE(_03630_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08347__B1 (.DIODE(_03628_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__A2 (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA__08348__B2 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08349__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08350__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08351__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08352__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08353__A2 (.DIODE(_03636_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A1 (.DIODE(\u_glbl_reg.reg_rdata[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08354__B1 (.DIODE(net1785));
 sky130_fd_sc_hd__diode_2 ANTENNA__08355__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08356__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08357__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08358__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08359__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08360__A2 (.DIODE(_03642_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__A2 (.DIODE(net584));
 sky130_fd_sc_hd__diode_2 ANTENNA__08361__B1 (.DIODE(_03640_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08362__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08363__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08364__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08365__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A1 (.DIODE(\u_gpio.reg_rdata[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08366__C1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08367__A2 (.DIODE(_03648_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08368__B1 (.DIODE(_03646_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08369__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08370__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08371__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08372__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A1 (.DIODE(\u_gpio.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08373__C1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A2 (.DIODE(_03654_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08374__A3 (.DIODE(_03655_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A1 (.DIODE(\u_glbl_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08375__B1 (.DIODE(net1781));
 sky130_fd_sc_hd__diode_2 ANTENNA__08376__A1 (.DIODE(net1088));
 sky130_fd_sc_hd__diode_2 ANTENNA__08377__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08378__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08379__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__A1 (.DIODE(\u_gpio.reg_rdata[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08380__C1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08381__A2 (.DIODE(_03660_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__A1 (.DIODE(net1798));
 sky130_fd_sc_hd__diode_2 ANTENNA__08382__B1 (.DIODE(_03658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08384__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08385__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08386__B (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A1 (.DIODE(\u_gpio.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08387__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08388__A2 (.DIODE(_03666_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__A1 (.DIODE(\u_glbl_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08389__B1 (.DIODE(net1808));
 sky130_fd_sc_hd__diode_2 ANTENNA__08391__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08392__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08393__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A1 (.DIODE(\u_gpio.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__A2 (.DIODE(net546));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08394__C1 (.DIODE(net541));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A1 (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA__08395__A2 (.DIODE(_03672_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08396__B1 (.DIODE(_03670_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08398__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08399__B2 (.DIODE(_03677_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08400__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A1 (.DIODE(\u_gpio.reg_rdata[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08401__C1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08402__A3 (.DIODE(_03679_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A1 (.DIODE(\u_glbl_reg.reg_rdata[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08403__B1 (.DIODE(net1777));
 sky130_fd_sc_hd__diode_2 ANTENNA__08405__B (.DIODE(net1207));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__A2 (.DIODE(net1119));
 sky130_fd_sc_hd__diode_2 ANTENNA__08406__B1 (.DIODE(net1114));
 sky130_fd_sc_hd__diode_2 ANTENNA__08407__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08408__C1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08409__A3 (.DIODE(_03685_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A1 (.DIODE(\u_glbl_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08410__B1 (.DIODE(_03682_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08412__B (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__A2 (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA__08413__B1 (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA__08414__B (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__A2 (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__B1 (.DIODE(net539));
 sky130_fd_sc_hd__diode_2 ANTENNA__08415__C1 (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA__08416__A3 (.DIODE(_03691_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__A2 (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA__08417__B1 (.DIODE(_03688_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08418__B (.DIODE(net1210));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__A2 (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA__08419__B1 (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA__08420__A2 (.DIODE(net1111));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A1 (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__A2 (.DIODE(net1110));
 sky130_fd_sc_hd__diode_2 ANTENNA__08421__B1 (.DIODE(net1091));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A1 (.DIODE(\u_timer.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08422__A2 (.DIODE(net723));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A1 (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__A2 (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA__08423__B1 (.DIODE(net553));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__A2 (.DIODE(_03471_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__B2 (.DIODE(net559));
 sky130_fd_sc_hd__diode_2 ANTENNA__08424__C1 (.DIODE(_03699_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__A (.DIODE(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08425__B (.DIODE(net548));
 sky130_fd_sc_hd__diode_2 ANTENNA__08426__A2 (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA__08427__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08449__B (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08450__A1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08455__B (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08457__A1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08460__B1 (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08461__A (.DIODE(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08473__A (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08474__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08475__S (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08476__S (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08477__S (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08478__S (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08479__S (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08480__S (.DIODE(_01198_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08481__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08483__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08485__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08487__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__A1 (.DIODE(_03408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08489__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08495__S (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08501__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08503__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08505__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08507__S (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA__08515__A1 (.DIODE(_03448_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08519__A0 (.DIODE(\u_ws281x.u_txd_0.led_data[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__A1 (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA__08521__B1 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08522__A2 (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08524__C (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA__08525__A (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08530__A1 (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08533__A1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08555__B (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08556__A1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08561__B (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08563__A1 (.DIODE(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08581__B (.DIODE(_03377_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__A1 (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08582__B1 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__A1 (.DIODE(_03382_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08583__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08584__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__A1 (.DIODE(_03388_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08585__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08586__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08587__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08588__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08589__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08590__S (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08591__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__A1 (.DIODE(_03402_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08593__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__A1 (.DIODE(_03405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08595__S (.DIODE(net731));
 sky130_fd_sc_hd__diode_2 ANTENNA__08613__A1 (.DIODE(_03432_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08615__A1 (.DIODE(_03435_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08617__A1 (.DIODE(_03440_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08621__A1 (.DIODE(_03445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08629__A1 (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08630__A2 (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08632__C (.DIODE(net570));
 sky130_fd_sc_hd__diode_2 ANTENNA__08633__A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08649__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08665__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08667__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08670__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08673__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08675__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08678__S (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08680__C_N (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08681__A2 (.DIODE(net521));
 sky130_fd_sc_hd__diode_2 ANTENNA__08703__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08706__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08708__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08711__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08714__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08716__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08719__S (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08721__C_N (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08722__A2 (.DIODE(net519));
 sky130_fd_sc_hd__diode_2 ANTENNA__08741__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08744__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08749__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08752__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08755__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08757__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08760__S (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08762__C_N (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08763__A2 (.DIODE(net515));
 sky130_fd_sc_hd__diode_2 ANTENNA__08845__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08846__A (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__S0 (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__08847__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08848__S (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__08849__S (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08850__A (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__A2 (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08851__B1 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08852__S (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__S0 (.DIODE(net1365));
 sky130_fd_sc_hd__diode_2 ANTENNA__08853__S1 (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA__08855__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08857__S (.DIODE(net1369));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__08858__B2 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08861__S (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08862__S (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__08865__S (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__A2 (.DIODE(net1226));
 sky130_fd_sc_hd__diode_2 ANTENNA__08867__B1 (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__A2 (.DIODE(_00999_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08868__B2 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__A1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__08869__B2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__A1 (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA__08871__C1 (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08872__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08873__S (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__08874__A (.DIODE(net1358));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__A1 (.DIODE(net1276));
 sky130_fd_sc_hd__diode_2 ANTENNA__08875__C1 (.DIODE(net1214));
 sky130_fd_sc_hd__diode_2 ANTENNA__08876__S1 (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08877__B2 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08878__A1 (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__08879__S (.DIODE(net1280));
 sky130_fd_sc_hd__diode_2 ANTENNA__08880__A2 (.DIODE(net1248));
 sky130_fd_sc_hd__diode_2 ANTENNA__08880__B1_N (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__08881__A (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__08882__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__08883__A (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__08884__A1 (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08885__S (.DIODE(net1275));
 sky130_fd_sc_hd__diode_2 ANTENNA__08886__B2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08889__A1 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08891__A1 (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA__08892__B2 (.DIODE(net1181));
 sky130_fd_sc_hd__diode_2 ANTENNA__08895__B2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__A2 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__08898__B2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__08900__B2 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08901__B2 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08902__B2 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08903__A1 (.DIODE(_00779_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08907__A1 (.DIODE(net1134));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__A (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA__08908__B (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08910__B1 (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A1 (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__08911__A2 (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08914__B1 (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A1 (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__08915__A2 (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08916__B (.DIODE(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08917__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_run ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08918__A (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A1 (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__08919__A2 (.DIODE(_03997_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__A (.DIODE(_01386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08920__B (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__A (.DIODE(_00873_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__B (.DIODE(_01386_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08921__C (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08926__A (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08938__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__A2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08942__B1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08944__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08946__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08947__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__A2 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08948__B1 (.DIODE(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08970__B (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08971__B1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08975__B (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08977__B1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08980__B1 (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08982__B1_N (.DIODE(net677));
 sky130_fd_sc_hd__diode_2 ANTENNA__08984__B (.DIODE(_01482_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__A (.DIODE(_00893_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08985__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08986__B (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08987__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08988__A (.DIODE(_00891_));
 sky130_fd_sc_hd__diode_2 ANTENNA__08989__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08990__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08991__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08992__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__08993__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08994__A (.DIODE(net726));
 sky130_fd_sc_hd__diode_2 ANTENNA__08995__B (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA__08996__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09000__A (.DIODE(_00885_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09002__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09004__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09006__A (.DIODE(_00882_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09010__A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09012__A (.DIODE(_00879_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09013__A_N (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09014__A1 (.DIODE(net1074));
 sky130_fd_sc_hd__diode_2 ANTENNA__09014__A2 (.DIODE(_01405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09016__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09018__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09030__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09034__B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09035__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09039__B (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09041__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09044__B1 (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09046__B1_N (.DIODE(net674));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__A_N (.DIODE(_01460_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09048__B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09049__A (.DIODE(_00913_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09052__A (.DIODE(net725));
 sky130_fd_sc_hd__diode_2 ANTENNA__09066__A1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09070__A2 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09072__A1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09074__A1 (.DIODE(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09076__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__09077__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__09078__A1 (.DIODE(net1072));
 sky130_fd_sc_hd__diode_2 ANTENNA__09080__B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09081__B1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09083__B1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09086__C (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09087__B1 (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09090__C (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09091__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09094__C (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09095__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09099__B (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09100__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09104__B (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA__09106__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09109__B1 (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09111__B1_N (.DIODE(net672));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09113__B (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09114__B (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09115__B (.DIODE(net1417));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09116__B (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__A (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09117__C_N (.DIODE(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09118__B (.DIODE(\u_gpio.cfg_gpio_dir_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09119__B (.DIODE(\u_gpio.cfg_gpio_dir_sel[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09120__B1_N (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09121__B1_N (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09122__B1_N (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09123__B1_N (.DIODE(\u_glbl_reg.cfg_multi_func_sel[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09124__B (.DIODE(net1406));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09125__B (.DIODE(net1408));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09126__B (.DIODE(net1410));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__09127__B (.DIODE(net1412));
 sky130_fd_sc_hd__diode_2 ANTENNA__09128__A1 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09129__D_N (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09130__B (.DIODE(net1651));
 sky130_fd_sc_hd__diode_2 ANTENNA__09131__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09132__B (.DIODE(_04107_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09133__D (.DIODE(\u_glbl_reg.cfg_multi_func_sel[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09134__B (.DIODE(_04108_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A1 (.DIODE(\u_gpio.cfg_gpio_dir_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A2 (.DIODE(\u_gpio.cfg_gpio_out_type[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09136__A3 (.DIODE(\u_glbl_reg.cfg_multi_func_sel[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__C (.DIODE(\u_glbl_reg.cfg_multi_func_sel[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09137__D (.DIODE(\u_glbl_reg.cfg_multi_func_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09138__B (.DIODE(_04109_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09139__C (.DIODE(\u_glbl_reg.cfg_multi_func_sel[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09140__B (.DIODE(_04110_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09142__B (.DIODE(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09143__B (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09144__B (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09145__B (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__A (.DIODE(net1109));
 sky130_fd_sc_hd__diode_2 ANTENNA__09146__B (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09148__A1 (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA__09151__B (.DIODE(\u_glbl_reg.u_random.s0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09152__B (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09157__B (.DIODE(\u_glbl_reg.u_random.s0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09162__B (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09186__B (.DIODE(\u_glbl_reg.u_random.s0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09191__A (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__A (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__09192__C (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__09196__A (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09206__A (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09213__B (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09219__A (.DIODE(\u_glbl_reg.u_random.s0[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09229__A (.DIODE(\u_glbl_reg.u_random.s0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09232__A (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09235__A (.DIODE(\u_glbl_reg.u_random.s0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09240__B (.DIODE(\u_glbl_reg.reg_3[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09241__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09242__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09245__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09246__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09247__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09251__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09252__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09253__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09255__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09256__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09257__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09258__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09259__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09260__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09261__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09262__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09263__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09264__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09265__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09266__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09267__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09268__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09269__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09270__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09271__A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__A (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09275__B (.DIODE(\u_glbl_reg.u_random.n1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__A (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09276__B (.DIODE(\u_glbl_reg.u_random.n1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__A (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09277__B (.DIODE(\u_glbl_reg.u_random.n1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__A (.DIODE(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09285__B (.DIODE(\u_glbl_reg.u_random.n1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__A (.DIODE(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09286__B (.DIODE(\u_glbl_reg.u_random.n1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__A (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09290__B (.DIODE(\u_glbl_reg.u_random.n1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__A (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09291__B (.DIODE(\u_glbl_reg.u_random.n1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__A (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09296__B (.DIODE(\u_glbl_reg.u_random.n1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__A (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09297__B (.DIODE(\u_glbl_reg.u_random.n1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__A (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09301__B (.DIODE(\u_glbl_reg.u_random.n1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__A (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09302__B (.DIODE(\u_glbl_reg.u_random.n1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__A (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09306__B (.DIODE(\u_glbl_reg.u_random.n1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09309__A (.DIODE(\u_glbl_reg.u_random.n0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09310__A (.DIODE(\u_glbl_reg.u_random.n0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A1 (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__A2 (.DIODE(\u_glbl_reg.u_random.n1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__B1 (.DIODE(\u_glbl_reg.u_random.n1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09312__C1 (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A1 (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09313__A2 (.DIODE(\u_glbl_reg.u_random.n1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09316__A (.DIODE(\u_glbl_reg.u_random.n0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09318__A (.DIODE(\u_glbl_reg.u_random.n0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__A (.DIODE(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09322__B (.DIODE(\u_glbl_reg.u_random.n1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__A (.DIODE(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09323__B (.DIODE(\u_glbl_reg.u_random.n1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09327__A (.DIODE(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09328__A (.DIODE(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__A (.DIODE(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09332__B (.DIODE(\u_glbl_reg.u_random.n1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__A (.DIODE(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09333__B (.DIODE(\u_glbl_reg.u_random.n1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__A (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09342__B (.DIODE(\u_glbl_reg.u_random.n1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__A (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09343__B (.DIODE(\u_glbl_reg.u_random.n1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__A (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09344__B (.DIODE(\u_glbl_reg.u_random.n1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__A (.DIODE(\u_glbl_reg.u_random.n0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09348__B (.DIODE(\u_glbl_reg.u_random.n1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__A (.DIODE(\u_glbl_reg.u_random.n0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09349__B (.DIODE(\u_glbl_reg.u_random.n1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__A (.DIODE(\u_glbl_reg.u_random.n0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09365__B (.DIODE(\u_glbl_reg.u_random.n1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__A (.DIODE(\u_glbl_reg.u_random.n0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09366__B (.DIODE(\u_glbl_reg.u_random.n1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09368__A (.DIODE(_04210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09369__A (.DIODE(\u_glbl_reg.u_random.n0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09371__A (.DIODE(\u_glbl_reg.u_random.n0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09373__A1 (.DIODE(_04210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__A (.DIODE(\u_glbl_reg.u_random.n0[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09375__B (.DIODE(\u_glbl_reg.u_random.n1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__A (.DIODE(\u_glbl_reg.u_random.n0[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09376__B (.DIODE(\u_glbl_reg.u_random.n1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__A (.DIODE(\u_glbl_reg.u_random.n0[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09377__B (.DIODE(\u_glbl_reg.u_random.n1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09380__A (.DIODE(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09383__A (.DIODE(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09384__A (.DIODE(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09388__A1 (.DIODE(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09389__A1 (.DIODE(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09391__A1 (.DIODE(_04210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09393__A (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09394__A (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09395__A (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09399__A (.DIODE(\u_glbl_reg.u_random.n0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09400__A (.DIODE(\u_glbl_reg.u_random.n0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09406__A (.DIODE(\u_glbl_reg.u_random.n0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09407__A (.DIODE(\u_glbl_reg.u_random.n0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09416__A1 (.DIODE(_04210_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__A (.DIODE(\u_glbl_reg.u_random.n0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09417__B (.DIODE(\u_glbl_reg.u_random.n1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__A (.DIODE(\u_glbl_reg.u_random.n0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09418__B (.DIODE(\u_glbl_reg.u_random.n1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__A (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09421__B (.DIODE(\u_glbl_reg.u_random.n1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__A (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09422__B (.DIODE(\u_glbl_reg.u_random.n1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__A (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09423__B (.DIODE(\u_glbl_reg.u_random.n1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__A (.DIODE(\u_glbl_reg.u_random.n0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09427__B (.DIODE(\u_glbl_reg.u_random.n1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__A (.DIODE(\u_glbl_reg.u_random.n0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09428__B (.DIODE(\u_glbl_reg.u_random.n1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__A (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09446__B (.DIODE(\u_glbl_reg.u_random.n1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__A (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09447__B (.DIODE(\u_glbl_reg.u_random.n1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09451__A (.DIODE(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09452__A (.DIODE(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09457__A (.DIODE(\u_glbl_reg.u_random.n0[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09458__B (.DIODE(_04288_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__A (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__09459__B (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A2 (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__A3 (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09460__B1 (.DIODE(_01559_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__A1 (.DIODE(_00850_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__A2 (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__A3 (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09461__B1 (.DIODE(_00776_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__B (.DIODE(_01270_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09463__C (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09464__A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09465__B (.DIODE(_00589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09466__B (.DIODE(_00589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09467__A (.DIODE(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__B (.DIODE(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__C (.DIODE(net1158));
 sky130_fd_sc_hd__diode_2 ANTENNA__09470__D (.DIODE(_01390_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09471__B (.DIODE(_01040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09472__A2 (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09473__A3 (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A0 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A1 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A2 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09474__A3 (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09478__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09479__A (.DIODE(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09480__B (.DIODE(_01040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09481__A2 (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09482__A3 (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A0 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A1 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A2 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09483__A3 (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09487__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09488__A (.DIODE(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09489__B (.DIODE(_01040_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__A2 (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09490__B1_N (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A2 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09491__A3 (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A0 (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A1 (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A2 (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__A3 (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S0 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09492__S1 (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A0 (.DIODE(_04308_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09493__A1 (.DIODE(_04307_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09494__B1 (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09495__B1 (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09496__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09497__C (.DIODE(_04309_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09498__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09499__B (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09500__B2 (.DIODE(net1135));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09502__B (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09503__B2 (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09505__B (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09506__B2 (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09508__B (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A1 (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA__09509__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09511__C (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A1 (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09512__A2 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__09513__B1 (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09514__B (.DIODE(_01001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09515__A1 (.DIODE(_01001_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09517__B (.DIODE(net666));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B1 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09518__B2 (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__A (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__C (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09520__D (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A1 (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A2 (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA__09521__A3 (.DIODE(net1145));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A1 (.DIODE(net670));
 sky130_fd_sc_hd__diode_2 ANTENNA__09522__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__A (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__09523__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__A (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__09524__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__A (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__09525__B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__A (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__09526__B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__A (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__09527__B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__09528__A (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__A (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__09529__B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__09530__A (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__09531__A (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__09532__A (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__A (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__09533__B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__A (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__09534__B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__09535__A (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__A (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__09536__B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09537__A (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__A (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__09538__B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__A (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__09539__B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__09540__A (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__09541__A (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__A (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__09542__B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09543__B (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A1 (.DIODE(net662));
 sky130_fd_sc_hd__diode_2 ANTENNA__09544__A2 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09546__C (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A1 (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09547__A2 (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A1 (.DIODE(net1179));
 sky130_fd_sc_hd__diode_2 ANTENNA__09548__A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09549__C (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A1 (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09550__A2 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A1 (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__09551__A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09552__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09554__A3 (.DIODE(net579));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__B (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09555__C (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A1 (.DIODE(net1249));
 sky130_fd_sc_hd__diode_2 ANTENNA__09557__A2 (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__A (.DIODE(net1299));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__B (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09558__C (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A1 (.DIODE(net1180));
 sky130_fd_sc_hd__diode_2 ANTENNA__09560__A2 (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__B (.DIODE(net1160));
 sky130_fd_sc_hd__diode_2 ANTENNA__09561__C (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A1 (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA__09563__A2 (.DIODE(_01144_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09564__A (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__09565__A (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__09566__A (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__09567__A (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__09568__A (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__09572__D (.DIODE(net1346));
 sky130_fd_sc_hd__diode_2 ANTENNA__09573__D (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__09574__D (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__09591__D (.DIODE(\u_gpio.u_bit[0].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09595__D (.DIODE(\u_gpio.u_bit[4].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09598__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09600__RESET_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__09604__D (.DIODE(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09605__D (.DIODE(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09606__D (.DIODE(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09608__D (.DIODE(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09609__D (.DIODE(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09610__D (.DIODE(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09612__D (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09614__D (.DIODE(\u_gpio.u_bit[27].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09615__D (.DIODE(\u_gpio.u_bit[28].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA__09617__RESET_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__09619__D (.DIODE(net1392));
 sky130_fd_sc_hd__diode_2 ANTENNA__09623__D (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__09627__D (.DIODE(net1417));
 sky130_fd_sc_hd__diode_2 ANTENNA__09631__D (.DIODE(net1403));
 sky130_fd_sc_hd__diode_2 ANTENNA__09635__D (.DIODE(net1400));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__D (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__09639__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__09643__D (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__D (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA__09647__RESET_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA__09651__D (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA__09655__D (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA__09659__D (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA__09663__D (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA__09667__D (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__D (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA__09671__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__09672__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__09673__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__09675__D (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA__09679__D (.DIODE(net1388));
 sky130_fd_sc_hd__diode_2 ANTENNA__09683__D (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA__09687__D (.DIODE(net1387));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__D (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA__09691__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__D (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA__09695__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09696__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09697__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09698__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09699__D (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA__09703__D (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA__09707__D (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__09710__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__09711__D (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__09715__D (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA__09719__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09720__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__09723__D (.DIODE(net1650));
 sky130_fd_sc_hd__diode_2 ANTENNA__09727__D (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__09732__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09733__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09734__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09735__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09736__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09737__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09738__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09739__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09740__RESET_B (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA__09741__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09742__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09743__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09744__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09745__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09746__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__09747__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09748__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09749__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09750__RESET_B (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA__09751__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09752__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09753__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09754__CLK (.DIODE(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09755__CLK (.DIODE(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09762__CLK (.DIODE(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__CLK (.DIODE(clknet_1_0__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09764__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__CLK (.DIODE(clknet_1_1__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09765__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__CLK (.DIODE(clknet_1_0__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09766__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__CLK (.DIODE(clknet_1_1__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09767__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__09768__CLK (.DIODE(clknet_1_0__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__CLK (.DIODE(clknet_1_1__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09769__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__09770__CLK (.DIODE(clknet_1_0__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__CLK (.DIODE(clknet_1_1__leaf__04546_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09771__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__09772__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__09773__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__09774__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__09775__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09776__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09777__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__09778__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09779__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__09780__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09781__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__09782__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09783__D (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09784__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__09785__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09786__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09787__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__09789__D (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09790__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09792__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09794__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09795__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__09796__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09797__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09798__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__09799__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__09801__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__09803__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__09804__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__09805__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__09806__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__09807__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09808__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__09809__RESET_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__09810__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__09811__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__09812__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09813__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__09814__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09815__D (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__09816__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09817__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__09818__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09819__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__09821__D (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__09822__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09824__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09826__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09827__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__09828__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09829__D (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__09830__D (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09831__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__09833__D (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__09834__D (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__09835__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__09836__D (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__D (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__09837__RESET_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__D (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__09838__RESET_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__09839__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__09840__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__09841__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__09842__D (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA__09843__D (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA__09844__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09845__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__09846__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09847__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09848__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__09849__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09850__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09851__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09853__D (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__09854__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09856__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09858__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09859__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__09861__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09869__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__09875__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__09876__RESET_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__09881__RESET_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__09892__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09893__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__09894__D (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09895__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__09897__D (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__09899__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__09900__D (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__09901__D (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__09902__D (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__09903__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09904__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__09905__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__09906__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__09907__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__09908__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09909__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__09910__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09911__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09912__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__09913__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09914__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09915__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09917__D (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09918__RESET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__09919__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09920__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09922__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09923__D (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09924__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__09925__D (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__D (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09926__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__09927__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__09929__D (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__09931__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__09932__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__09933__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__09934__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__09935__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09936__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__09937__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__09938__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__09939__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__09940__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09941__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09942__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__09943__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09944__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__09945__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09946__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09947__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__CLK (.DIODE(clknet_1_0__leaf__04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09949__D (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__CLK (.DIODE(clknet_1_0__leaf__04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09950__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__CLK (.DIODE(clknet_1_0__leaf__04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09951__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09952__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09953__CLK (.DIODE(clknet_1_0__leaf__04501_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09954__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__D (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09955__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__09956__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__D (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__09957__RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__D (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__09958__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__09959__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__09961__D (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__09962__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__09963__D (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA__09964__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__09965__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__09966__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__09967__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__09968__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__09969__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__09970__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__09971__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__09972__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__09973__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__09974__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__09975__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__09976__D (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__09977__RESET_B (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA__09978__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__09979__RESET_B (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__CLK (.DIODE(clknet_1_0__leaf__04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09981__D (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__CLK (.DIODE(clknet_1_0__leaf__04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__D (.DIODE(net1287));
 sky130_fd_sc_hd__diode_2 ANTENNA__09982__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__CLK (.DIODE(clknet_1_0__leaf__04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__09983__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__09984__D (.DIODE(net1637));
 sky130_fd_sc_hd__diode_2 ANTENNA__09985__CLK (.DIODE(clknet_1_0__leaf__04497_));
 sky130_fd_sc_hd__diode_2 ANTENNA__09986__D (.DIODE(net1622));
 sky130_fd_sc_hd__diode_2 ANTENNA__09987__D (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__09988__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09989__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09990__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09991__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09992__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09993__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09994__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09995__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09996__RESET_B (.DIODE(net1386));
 sky130_fd_sc_hd__diode_2 ANTENNA__09997__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__09998__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__09999__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10000__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10001__RESET_B (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10002__RESET_B (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10003__RESET_B (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10004__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10005__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10007__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__10008__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__10009__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__10010__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__10011__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10012__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10013__RESET_B (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA__10014__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10015__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10016__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10017__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10018__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10025__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10026__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10028__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10029__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10030__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10031__RESET_B (.DIODE(net913));
 sky130_fd_sc_hd__diode_2 ANTENNA__10032__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10033__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10034__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10035__RESET_B (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10036__D (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10046__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10050__D (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10055__D (.DIODE(\u_glbl_reg.u_random.s1_xor_s0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10061__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10080__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10090__RESET_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__10091__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10097__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10100__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10101__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10102__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10103__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10104__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10105__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10106__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10107__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10108__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10109__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10110__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10111__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10112__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10113__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10114__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10115__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10116__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10117__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10118__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10119__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10120__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10121__CLK (.DIODE(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10122__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10123__CLK (.DIODE(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10124__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10125__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10126__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10127__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10128__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10129__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10130__CLK (.DIODE(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10131__CLK (.DIODE(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10132__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10133__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10134__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10135__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10136__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10137__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10138__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10139__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10140__D (.DIODE(net1889));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10141__D (.DIODE(net1881));
 sky130_fd_sc_hd__diode_2 ANTENNA__10142__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10143__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10144__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10145__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10146__D (.DIODE(net1909));
 sky130_fd_sc_hd__diode_2 ANTENNA__10147__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10148__D (.DIODE(net1917));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10149__D (.DIODE(net1884));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10150__D (.DIODE(net1931));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__D (.DIODE(net1927));
 sky130_fd_sc_hd__diode_2 ANTENNA__10151__RESET_B (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA__10152__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10153__CLK (.DIODE(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10154__D (.DIODE(net1928));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__CLK (.DIODE(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10155__D (.DIODE(net1905));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10156__D (.DIODE(net1892));
 sky130_fd_sc_hd__diode_2 ANTENNA__10157__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__D (.DIODE(net1915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10158__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10159__D (.DIODE(net1894));
 sky130_fd_sc_hd__diode_2 ANTENNA__10160__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10161__RESET_B (.DIODE(net947));
 sky130_fd_sc_hd__diode_2 ANTENNA__10162__CLK (.DIODE(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10163__CLK (.DIODE(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10166__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10167__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10176__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10177__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__10179__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__10184__RESET_B (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA__10189__RESET_B (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA__10193__CLK (.DIODE(clknet_1_0__leaf__04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10194__CLK (.DIODE(clknet_1_0__leaf__04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__CLK (.DIODE(clknet_1_0__leaf__04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10195__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10196__CLK (.DIODE(clknet_1_0__leaf__04395_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10199__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10200__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10201__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10203__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10205__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10211__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10212__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10213__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10214__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10223__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10224__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10225__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10226__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10227__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10228__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10229__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10230__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10231__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10232__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10233__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10234__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10235__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10236__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10237__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10238__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10239__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10240__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10241__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10242__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10243__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10244__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10245__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10246__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10247__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10248__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10249__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10250__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10251__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10252__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10253__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10254__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__CLK (.DIODE(clknet_1_0__leaf__04403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__D (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10255__RESET_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__10256__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__CLK (.DIODE(clknet_1_0__leaf__04403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10258__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__CLK (.DIODE(clknet_1_0__leaf__04403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10259__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10260__D (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__CLK (.DIODE(clknet_1_0__leaf__04403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10261__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10262__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__10263__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10264__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10265__SET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10266__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10267__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10268__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10269__SET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10270__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10271__RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10272__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10273__SET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10274__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10275__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10276__RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10277__SET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10278__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10279__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10280__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10281__D (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10282__RESET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10283__SET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10284__SET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10285__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10286__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10287__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10288__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10289__RESET_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10290__RESET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10291__RESET_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10292__SET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10293__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10294__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__CLK (.DIODE(clknet_1_0__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10295__D (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__CLK (.DIODE(clknet_1_1__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10296__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__CLK (.DIODE(clknet_1_1__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10297__RESET_B (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__CLK (.DIODE(clknet_1_0__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10298__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__CLK (.DIODE(clknet_1_1__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10299__RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__CLK (.DIODE(clknet_1_0__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10300__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__CLK (.DIODE(clknet_1_1__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10301__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__CLK (.DIODE(clknet_1_0__leaf__04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10302__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10303__RESET_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__CLK (.DIODE(clknet_1_1__leaf__04405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10304__RESET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__10305__CLK (.DIODE(clknet_1_1__leaf__04405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10306__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10307__SET_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__CLK (.DIODE(clknet_1_1__leaf__04405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10308__D (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__CLK (.DIODE(clknet_1_1__leaf__04405_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10309__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10310__RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10311__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10312__SET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10313__SET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10314__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10315__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10316__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10317__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__10318__RESET_B (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10319__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10320__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10321__RESET_B (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA__10322__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10323__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10324__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10325__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10326__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__CLK (.DIODE(clknet_1_1__leaf__04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10327__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__D (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10328__SET_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__CLK (.DIODE(clknet_1_1__leaf__04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10329__SET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__CLK (.DIODE(clknet_1_1__leaf__04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10330__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10331__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10332__RESET_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__CLK (.DIODE(clknet_1_1__leaf__04410_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10333__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10334__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10335__RESET_B (.DIODE(net1044));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10336__RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10337__RESET_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10338__RESET_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10339__RESET_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10340__RESET_B (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10341__RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10342__RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__CLK (.DIODE(clknet_1_1__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10343__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__CLK (.DIODE(clknet_1_0__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10344__D (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__CLK (.DIODE(clknet_1_1__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10345__RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__CLK (.DIODE(clknet_1_0__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10346__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__CLK (.DIODE(clknet_1_1__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10347__SET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__CLK (.DIODE(clknet_1_0__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10348__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__CLK (.DIODE(clknet_1_1__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10349__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__CLK (.DIODE(clknet_1_0__leaf__04408_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10350__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10351__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10352__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10353__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10354__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10355__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10356__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10357__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__D (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__10358__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__CLK (.DIODE(clknet_1_0__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10359__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__CLK (.DIODE(clknet_1_1__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10360__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__CLK (.DIODE(clknet_1_0__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10361__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__CLK (.DIODE(clknet_1_1__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10362__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__CLK (.DIODE(clknet_1_0__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10363__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__CLK (.DIODE(clknet_1_0__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10364__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__CLK (.DIODE(clknet_1_1__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10365__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__CLK (.DIODE(clknet_1_1__leaf__04414_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10366__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__D (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10367__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10368__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10369__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10370__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10371__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10372__D (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__10373__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10374__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__CLK (.DIODE(clknet_1_0__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10375__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__CLK (.DIODE(clknet_1_1__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10376__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__CLK (.DIODE(clknet_1_1__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10377__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__CLK (.DIODE(clknet_1_0__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10378__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__CLK (.DIODE(clknet_1_1__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10379__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__CLK (.DIODE(clknet_1_0__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10380__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__CLK (.DIODE(clknet_1_0__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10381__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__CLK (.DIODE(clknet_1_1__leaf__04412_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__10382__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__10403__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10404__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10405__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10406__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10407__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10408__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10409__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10410__RESET_B (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA__10411__RESET_B (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA__10412__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__10413__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10414__D (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10415__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10417__RESET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__10418__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10419__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10420__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10421__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10422__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10423__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10424__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10425__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10426__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__10427__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10428__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10429__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10430__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10431__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10432__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10433__D (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10434__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__10435__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10436__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10437__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10438__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10439__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10440__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10441__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10442__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10443__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10444__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__10445__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10446__D (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10447__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10449__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10450__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10451__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10452__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10453__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10454__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10455__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10456__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10457__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10458__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10459__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10460__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10461__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10462__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10463__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10464__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__D (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10465__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10466__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10467__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10468__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10469__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10470__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10471__D (.DIODE(net1636));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10472__RESET_B (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA__10473__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10474__D (.DIODE(net1615));
 sky130_fd_sc_hd__diode_2 ANTENNA__10475__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10476__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__D (.DIODE(net1488));
 sky130_fd_sc_hd__diode_2 ANTENNA__10477__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10478__D (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10479__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10481__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10482__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10483__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10484__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__CLK (.DIODE(clknet_1_1__leaf__04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10485__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__CLK (.DIODE(clknet_1_1__leaf__04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10486__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10487__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__CLK (.DIODE(clknet_1_1__leaf__04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__D (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__10488__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__CLK (.DIODE(clknet_1_1__leaf__04429_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10489__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10490__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10491__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10492__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__D (.DIODE(net1589));
 sky130_fd_sc_hd__diode_2 ANTENNA__10493__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10494__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10495__RESET_B (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA__10496__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__10497__D (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10498__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__10499__D (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__10500__D (.DIODE(net1418));
 sky130_fd_sc_hd__diode_2 ANTENNA__10501__D (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10502__RESET_B (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA__10503__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10504__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10505__D (.DIODE(net1621));
 sky130_fd_sc_hd__diode_2 ANTENNA__10506__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10508__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10509__D (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA__10510__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10511__RESET_B (.DIODE(net763));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10512__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10513__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10514__RESET_B (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10515__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10516__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10517__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10518__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10519__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10520__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10521__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10522__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10523__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__D (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10524__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10525__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10526__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10527__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10528__RESET_B (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10529__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10530__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10531__D (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__10532__D (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10533__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10534__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10535__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10536__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10537__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10538__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10539__D (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA__10540__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__10541__D (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__10542__D (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA__10543__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10545__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10546__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10547__D (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10548__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10549__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10550__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10551__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__10552__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10553__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10554__RESET_B (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10555__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10556__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10557__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__10558__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10559__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__D (.DIODE(net1556));
 sky130_fd_sc_hd__diode_2 ANTENNA__10560__RESET_B (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__D (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10561__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10562__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__D (.DIODE(net1534));
 sky130_fd_sc_hd__diode_2 ANTENNA__10563__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10564__RESET_B (.DIODE(net744));
 sky130_fd_sc_hd__diode_2 ANTENNA__10565__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10566__D (.DIODE(net1512));
 sky130_fd_sc_hd__diode_2 ANTENNA__10567__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10568__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10569__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10570__D (.DIODE(net1474));
 sky130_fd_sc_hd__diode_2 ANTENNA__10571__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__10572__D (.DIODE(net1598));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10573__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10574__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__D (.DIODE(net1566));
 sky130_fd_sc_hd__diode_2 ANTENNA__10575__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10576__D (.DIODE(net1559));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__D (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA__10577__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10578__D (.DIODE(net1545));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__D (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__10579__RESET_B (.DIODE(net777));
 sky130_fd_sc_hd__diode_2 ANTENNA__10580__D (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__10581__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10583__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10584__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10585__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10586__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10588__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__10589__D (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__D (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10590__RESET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__10591__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__D (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA__10592__RESET_B (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA__10593__D (.DIODE(net1442));
 sky130_fd_sc_hd__diode_2 ANTENNA__10594__D (.DIODE(net1434));
 sky130_fd_sc_hd__diode_2 ANTENNA__10595__D (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA__10596__D (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__10597__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10598__D (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA__10599__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10600__D (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA__10601__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10602__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__10603__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10604__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10605__D (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA__10606__D (.DIODE(net1466));
 sky130_fd_sc_hd__diode_2 ANTENNA__10607__D (.DIODE(net1457));
 sky130_fd_sc_hd__diode_2 ANTENNA__10608__D (.DIODE(net1448));
 sky130_fd_sc_hd__diode_2 ANTENNA__10609__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10610__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__CLK (.DIODE(clknet_1_1__leaf__04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__D (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10611__RESET_B (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__CLK (.DIODE(clknet_1_1__leaf__04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10612__D (.DIODE(net1526));
 sky130_fd_sc_hd__diode_2 ANTENNA__10613__D (.DIODE(net1519));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__CLK (.DIODE(clknet_1_1__leaf__04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10614__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10615__D (.DIODE(net1505));
 sky130_fd_sc_hd__diode_2 ANTENNA__10616__D (.DIODE(net1498));
 sky130_fd_sc_hd__diode_2 ANTENNA__10617__D (.DIODE(net1481));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__CLK (.DIODE(clknet_1_1__leaf__04445_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10618__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__D (.DIODE(net1603));
 sky130_fd_sc_hd__diode_2 ANTENNA__10619__RESET_B (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA__10620__D (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10621__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10622__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10623__RESET_B (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA__10624__D (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__10625__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10626__RESET_B (.DIODE(net898));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__D (.DIODE(net1293));
 sky130_fd_sc_hd__diode_2 ANTENNA__10627__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__D (.DIODE(net1572));
 sky130_fd_sc_hd__diode_2 ANTENNA__10628__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__D (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA__10629__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__CLK (.DIODE(clknet_1_1__leaf__04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__D (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA__10630__SET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__CLK (.DIODE(clknet_1_1__leaf__04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__D (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA__10631__RESET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__CLK (.DIODE(clknet_1_1__leaf__04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10632__RESET_B (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__D (.DIODE(net1441));
 sky130_fd_sc_hd__diode_2 ANTENNA__10633__RESET_B (.DIODE(net1046));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__CLK (.DIODE(clknet_1_1__leaf__04451_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10634__D (.DIODE(net1433));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__D (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA__10635__RESET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__D (.DIODE(net1527));
 sky130_fd_sc_hd__diode_2 ANTENNA__10636__RESET_B (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA__10638__D (.DIODE(net1513));
 sky130_fd_sc_hd__diode_2 ANTENNA__10639__D (.DIODE(net1506));
 sky130_fd_sc_hd__diode_2 ANTENNA__10640__D (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__D (.DIODE(net1482));
 sky130_fd_sc_hd__diode_2 ANTENNA__10641__RESET_B (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA__10642__D (.DIODE(net1475));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__D (.DIODE(net1604));
 sky130_fd_sc_hd__diode_2 ANTENNA__10643__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__D (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA__10644__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__D (.DIODE(net1586));
 sky130_fd_sc_hd__diode_2 ANTENNA__10645__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__D (.DIODE(net1579));
 sky130_fd_sc_hd__diode_2 ANTENNA__10646__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__10647__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__D (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA__10648__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__D (.DIODE(net1549));
 sky130_fd_sc_hd__diode_2 ANTENNA__10649__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__D (.DIODE(net1541));
 sky130_fd_sc_hd__diode_2 ANTENNA__10650__RESET_B (.DIODE(net1062));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__D (.DIODE(net1425));
 sky130_fd_sc_hd__diode_2 ANTENNA__10651__RESET_B (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__D (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA__10652__RESET_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__D (.DIODE(net1286));
 sky130_fd_sc_hd__diode_2 ANTENNA__10653__RESET_B (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__D (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA__10654__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10655__D (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__D (.DIODE(net1628));
 sky130_fd_sc_hd__diode_2 ANTENNA__10656__RESET_B (.DIODE(net1058));
 sky130_fd_sc_hd__diode_2 ANTENNA__10657__D (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__D (.DIODE(net1614));
 sky130_fd_sc_hd__diode_2 ANTENNA__10658__RESET_B (.DIODE(net1059));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10659__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__D (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__10660__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__10661__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__10662__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__10663__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__10664__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__10665__RESET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__10666__SET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10667__D (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__10668__D (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA__10669__D (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10670__D (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10671__D (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10672__D (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA__10673__D (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA__10674__D (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10675__SET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10676__RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10677__SET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10678__RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10679__SET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10680__RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10681__RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10682__RESET_B (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA__10683__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__10684__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__10685__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__10686__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__10687__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__D (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA__10688__SET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__10689__SET_B (.DIODE(net1064));
 sky130_fd_sc_hd__diode_2 ANTENNA__10690__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__10691__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10692__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10693__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10694__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10695__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10696__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10697__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10698__RESET_B (.DIODE(net752));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__D (.DIODE(net1306));
 sky130_fd_sc_hd__diode_2 ANTENNA__10702__GATE_N (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__D (.DIODE(net1305));
 sky130_fd_sc_hd__diode_2 ANTENNA__10703__GATE_N (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__D (.DIODE(net1304));
 sky130_fd_sc_hd__diode_2 ANTENNA__10704__GATE_N (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__D (.DIODE(net1650));
 sky130_fd_sc_hd__diode_2 ANTENNA__10705__GATE_N (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__D (.DIODE(net1571));
 sky130_fd_sc_hd__diode_2 ANTENNA__10706__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__D (.DIODE(net1497));
 sky130_fd_sc_hd__diode_2 ANTENNA__10707__GATE_N (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__D (.DIODE(net1417));
 sky130_fd_sc_hd__diode_2 ANTENNA__10708__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__D (.DIODE(net1403));
 sky130_fd_sc_hd__diode_2 ANTENNA__10709__GATE_N (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__D (.DIODE(net1397));
 sky130_fd_sc_hd__diode_2 ANTENNA__10710__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__D (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA__10711__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__D (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA__10712__GATE_N (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__D (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA__10713__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10714__D (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__D (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA__10715__GATE_N (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__D (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__10716__GATE_N (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__D (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA__10717__GATE_N (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA__10718__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10719__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10720__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10721__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10723__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10724__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10725__RESET_B (.DIODE(net1378));
 sky130_fd_sc_hd__diode_2 ANTENNA__10726__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10728__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10730__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10734__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10735__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10736__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10737__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10738__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10739__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10740__RESET_B (.DIODE(net1382));
 sky130_fd_sc_hd__diode_2 ANTENNA__10741__RESET_B (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA__10742__RESET_B (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10743__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10744__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10745__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10746__RESET_B (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA__10747__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10748__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10749__RESET_B (.DIODE(net1380));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__D (.DIODE(net2318));
 sky130_fd_sc_hd__diode_2 ANTENNA__10761__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10762__D (.DIODE(net2063));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10763__D (.DIODE(\u_glbl_reg.reg_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10764__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10765__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__D (.DIODE(\u_glbl_reg.reg_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10766__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10767__D (.DIODE(\u_glbl_reg.reg_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__CLK (.DIODE(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10768__D (.DIODE(\u_glbl_reg.reg_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10769__RESET_B (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10770__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10771__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10772__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10773__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10774__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10775__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10776__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10777__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10778__RESET_B (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA__10779__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10780__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10781__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10782__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10783__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10784__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10785__CLK (.DIODE(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10786__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10787__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10788__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__CLK (.DIODE(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10789__RESET_B (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA__10790__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10791__D (.DIODE(\u_glbl_reg.reg_out[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__CLK (.DIODE(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10792__D (.DIODE(\u_glbl_reg.reg_out[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10793__RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__D (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 ANTENNA__10798__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__10801__D (.DIODE(\u_glbl_reg.ir_intr_s ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10807__RESET_B (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA__10814__GATE (.DIODE(net1307));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__D (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__10815__RESET_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__D (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__10816__RESET_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__10817__D (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__D (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__10818__RESET_B (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA__10819__D (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__D (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10822__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__D (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10823__RESET_B (.DIODE(net902));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__D (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10824__RESET_B (.DIODE(net915));
 sky130_fd_sc_hd__diode_2 ANTENNA__10825__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__D (.DIODE(\u_ws281x.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10826__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__D (.DIODE(\u_ws281x.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10827__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__10828__D (.DIODE(\u_ws281x.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10829__D (.DIODE(\u_ws281x.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10830__D (.DIODE(\u_ws281x.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10831__D (.DIODE(\u_ws281x.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10832__D (.DIODE(\u_ws281x.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10833__D (.DIODE(\u_ws281x.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__10858__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10859__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10860__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__10861__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10862__D (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10863__D (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__10864__D (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10865__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__10866__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__10867__D (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__10868__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__10869__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__10870__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__10871__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__10872__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__10873__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__10874__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__10875__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__10876__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10877__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__10878__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10878__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__10879__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__10880__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__10881__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__10882__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10883__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10884__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10885__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10886__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10887__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10888__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10889__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10890__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10891__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10892__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__10893__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10894__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10895__RESET_B (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10896__RESET_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__10897__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10898__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__10899__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__10900__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10901__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__10902__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10903__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__10904__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__10905__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__10906__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__10907__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__10908__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__10909__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__10910__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__10911__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10914__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10915__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10916__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10917__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10918__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10919__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10920__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10921__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10922__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10923__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10924__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10925__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__CLK (.DIODE(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10926__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10927__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10928__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10929__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10930__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10931__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10932__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10933__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10934__D (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10935__D (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10936__D (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__CLK (.DIODE(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10937__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10938__D (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10939__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10940__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10941__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10942__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10943__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10944__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10945__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10946__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10947__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10948__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10949__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__CLK (.DIODE(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10950__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10951__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10952__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10953__D (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10954__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10955__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10956__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10957__D (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10958__D (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10959__D (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10960__D (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__CLK (.DIODE(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10961__D (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__10962__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__10963__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__10964__SET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__10965__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10966__D (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10967__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10968__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10969__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10970__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10971__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10972__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10973__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10974__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10975__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10976__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__CLK (.DIODE(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10977__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10978__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10979__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10980__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10981__D (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10982__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10983__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10984__D (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10985__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10986__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10987__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10988__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__CLK (.DIODE(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10989__D (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10990__D (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10991__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10992__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10993__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10994__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10995__D (.DIODE(net1455));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10996__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10997__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10998__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__10999__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11000__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11001__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11002__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11003__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11004__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11005__D (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11006__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11007__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11008__D (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11009__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11010__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11011__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__CLK (.DIODE(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11012__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__CLK (.DIODE(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11013__D (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__11015__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11016__RESET_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__11017__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11018__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11019__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11020__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11021__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11022__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__11023__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__11024__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__11025__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__11026__RESET_B (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA__11033__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11034__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11035__RESET_B (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA__11036__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11037__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11038__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11039__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11040__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11041__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11044__RESET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11045__RESET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11049__RESET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11050__RESET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11057__SET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11058__SET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11059__SET_B (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA__11065__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11066__RESET_B (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA__11067__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11068__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11069__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11070__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11071__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11072__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11073__RESET_B (.DIODE(net1029));
 sky130_fd_sc_hd__diode_2 ANTENNA__11074__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11075__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11076__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11077__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11078__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11079__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11081__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11085__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11086__RESET_B (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA__11087__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11088__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11089__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11099__RESET_B (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA__11130__RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__11131__RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__11140__RESET_B (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11142__D (.DIODE(\u_timer.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11143__D (.DIODE(\u_timer.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11144__D (.DIODE(\u_timer.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11145__D (.DIODE(\u_timer.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11146__D (.DIODE(\u_timer.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11147__D (.DIODE(\u_timer.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11148__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11149__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11150__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11151__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11152__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11153__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11154__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11155__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11156__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11157__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11158__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11159__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11160__RESET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__11161__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11162__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__CLK (.DIODE(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11163__RESET_B (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA__11164__CLK (.DIODE(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11165__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11166__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11167__RESET_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__11168__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11169__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11170__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11171__RESET_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__11172__CLK (.DIODE(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11173__CLK (.DIODE(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11174__D (.DIODE(net1606));
 sky130_fd_sc_hd__diode_2 ANTENNA__11175__D (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11176__D (.DIODE(net1590));
 sky130_fd_sc_hd__diode_2 ANTENNA__11177__D (.DIODE(net1581));
 sky130_fd_sc_hd__diode_2 ANTENNA__11178__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11179__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11180__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11181__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11182__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11183__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11184__D (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__11185__D (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__11186__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__11187__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11188__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11189__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11190__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__11191__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__11192__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__11193__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__11194__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__D (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA__11195__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__11196__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11197__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__11198__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11199__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11200__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11201__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__11202__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11203__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__11204__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__11205__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11206__D (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA__11207__D (.DIODE(net1599));
 sky130_fd_sc_hd__diode_2 ANTENNA__11208__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__D (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA__11209__RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__11210__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11211__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11212__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11213__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11214__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11215__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11216__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__11217__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11218__D (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__11219__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11220__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11221__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11222__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__11223__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__11224__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__11225__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__11226__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__D (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA__11227__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11228__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__11229__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__11230__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11231__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11232__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11233__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__11234__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11235__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__11236__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__11237__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11238__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11239__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__11240__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11241__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11242__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11243__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11244__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11245__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11246__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11247__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11248__D (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA__11249__D (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA__11250__D (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__11251__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11252__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11253__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11254__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__11255__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__11256__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__11257__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__11258__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__11259__D (.DIODE(net1455));
 sky130_fd_sc_hd__diode_2 ANTENNA__11260__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__11261__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__11262__D (.DIODE(net1431));
 sky130_fd_sc_hd__diode_2 ANTENNA__11263__D (.DIODE(net1424));
 sky130_fd_sc_hd__diode_2 ANTENNA__11264__D (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA__11265__D (.DIODE(net1649));
 sky130_fd_sc_hd__diode_2 ANTENNA__11266__D (.DIODE(net1640));
 sky130_fd_sc_hd__diode_2 ANTENNA__11267__D (.DIODE(net1634));
 sky130_fd_sc_hd__diode_2 ANTENNA__11268__D (.DIODE(net1625));
 sky130_fd_sc_hd__diode_2 ANTENNA__11269__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11270__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11271__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__11272__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11273__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11274__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11275__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11276__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11277__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11278__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11279__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11280__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__11281__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11282__D (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__D (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA__11283__RESET_B (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA__11284__D (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA__11285__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11286__D (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__11287__D (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__11288__D (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__11289__D (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__11290__D (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__11291__D (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA__11292__D (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__11293__D (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__11294__D (.DIODE(net1429));
 sky130_fd_sc_hd__diode_2 ANTENNA__11295__D (.DIODE(net1423));
 sky130_fd_sc_hd__diode_2 ANTENNA__11296__D (.DIODE(net1291));
 sky130_fd_sc_hd__diode_2 ANTENNA__11297__D (.DIODE(net1647));
 sky130_fd_sc_hd__diode_2 ANTENNA__11298__D (.DIODE(net1642));
 sky130_fd_sc_hd__diode_2 ANTENNA__11299__D (.DIODE(net1632));
 sky130_fd_sc_hd__diode_2 ANTENNA__11300__D (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA__11301__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11326__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11335__RESET_B (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA__11343__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11344__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11345__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11346__RESET_B (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA__11370__D (.DIODE(\u_semaphore.reg_out[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11378__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11381__RESET_B (.DIODE(net1018));
 sky130_fd_sc_hd__diode_2 ANTENNA__11384__CLK (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__11390__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11391__D (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__11392__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11393__D (.DIODE(net1296));
 sky130_fd_sc_hd__diode_2 ANTENNA__11394__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11395__D (.DIODE(net1490));
 sky130_fd_sc_hd__diode_2 ANTENNA__11396__D (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11397__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11398__D (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__11399__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11400__D (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__11401__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__11404__D (.DIODE(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11405__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11406__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11407__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11408__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11409__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11410__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11411__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11412__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11413__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11414__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11415__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11416__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11417__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11418__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11419__CLK (.DIODE(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11420__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11421__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11422__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11423__CLK (.DIODE(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11426__RESET_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__11427__RESET_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__11440__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11441__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11442__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11443__CLK (.DIODE(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11444__CLK (.DIODE(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11445__CLK (.DIODE(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11446__CLK (.DIODE(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11447__CLK (.DIODE(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11457__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11458__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11459__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11461__CLK (.DIODE(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11472__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11473__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11474__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11475__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11476__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11477__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11478__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11479__D (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__11480__D (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__11481__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__11482__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__11483__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11484__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__11485__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__11486__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__11487__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__11488__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11489__D (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA__11490__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11491__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__11492__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11493__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__11494__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__11495__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11496__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11497__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__11498__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11499__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11500__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11501__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11502__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11503__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11504__D (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11505__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11506__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11507__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11508__D (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA__11509__D (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA__11510__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11511__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11512__D (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__11513__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__11514__RESET_B (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA__11515__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11516__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__11517__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__11518__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__11519__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__11520__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11521__D (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__11522__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11523__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__11524__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11525__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__11526__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__11527__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11528__D (.DIODE(net1607));
 sky130_fd_sc_hd__diode_2 ANTENNA__11529__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__11530__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11531__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11532__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11533__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11534__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11535__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11536__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11537__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11538__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11539__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11540__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11541__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11542__D (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11543__D (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__11544__D (.DIODE(net1300));
 sky130_fd_sc_hd__diode_2 ANTENNA__11545__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__11546__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__11547__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11548__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__11549__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__11550__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__11551__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__11552__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__D (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__11553__RESET_B (.DIODE(net1021));
 sky130_fd_sc_hd__diode_2 ANTENNA__11554__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11555__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__11556__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11557__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__11558__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__11559__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11560__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11561__D (.DIODE(net1600));
 sky130_fd_sc_hd__diode_2 ANTENNA__11562__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11563__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11564__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11565__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11566__D (.DIODE(net1553));
 sky130_fd_sc_hd__diode_2 ANTENNA__11567__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11568__D (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11569__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11570__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11571__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11572__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11573__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11574__D (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA__11575__D (.DIODE(net1618));
 sky130_fd_sc_hd__diode_2 ANTENNA__11576__D (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA__11577__D (.DIODE(net1578));
 sky130_fd_sc_hd__diode_2 ANTENNA__11578__D (.DIODE(net1493));
 sky130_fd_sc_hd__diode_2 ANTENNA__11579__D (.DIODE(net1470));
 sky130_fd_sc_hd__diode_2 ANTENNA__11580__D (.DIODE(net1464));
 sky130_fd_sc_hd__diode_2 ANTENNA__11581__D (.DIODE(net1453));
 sky130_fd_sc_hd__diode_2 ANTENNA__11582__D (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA__11583__D (.DIODE(net1439));
 sky130_fd_sc_hd__diode_2 ANTENNA__11584__D (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__11585__D (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__11586__D (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__11587__D (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__11588__D (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__11589__D (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__11590__D (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__11591__D (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__11592__D (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__11593__D (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__11594__D (.DIODE(net1591));
 sky130_fd_sc_hd__diode_2 ANTENNA__11595__D (.DIODE(net1583));
 sky130_fd_sc_hd__diode_2 ANTENNA__11596__D (.DIODE(net1568));
 sky130_fd_sc_hd__diode_2 ANTENNA__11597__D (.DIODE(net1561));
 sky130_fd_sc_hd__diode_2 ANTENNA__11598__D (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__11599__D (.DIODE(net1546));
 sky130_fd_sc_hd__diode_2 ANTENNA__11600__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11601__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11602__D (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11603__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11604__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11605__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11606__CLK (.DIODE(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11607__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11608__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11609__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11610__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11611__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11615__CLK (.DIODE(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11624__D (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11626__D (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11630__D (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11633__RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__11634__RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__11635__RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__11636__RESET_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__11637__RESET_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__11638__RESET_B (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA__11664__RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__11665__RESET_B (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA__11668__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11669__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11670__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11671__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11672__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11673__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11674__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11675__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11676__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11677__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11678__CLK (.DIODE(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11679__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11680__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11681__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11682__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11683__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11684__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11685__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__CLK (.DIODE(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11686__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11703__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11704__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11705__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11706__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11707__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11708__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11709__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11710__CLK (.DIODE(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11715__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11719__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11720__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11721__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11722__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11724__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11725__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11726__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11727__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11729__D (.DIODE(net2127));
 sky130_fd_sc_hd__diode_2 ANTENNA__11730__D (.DIODE(net2113));
 sky130_fd_sc_hd__diode_2 ANTENNA__11731__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__D (.DIODE(net2105));
 sky130_fd_sc_hd__diode_2 ANTENNA__11732__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__CLK (.DIODE(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11733__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11735__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11736__D (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11737__D (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11738__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11739__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11740__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11741__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11742__D (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__11743__D (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11744__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11745__D (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__11746__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__11747__D (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA__11748__D (.DIODE(net1450));
 sky130_fd_sc_hd__diode_2 ANTENNA__11749__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__11750__D (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11751__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11752__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11753__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__11754__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11755__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__11756__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11757__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11758__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11759__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11760__D (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__11761__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11762__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11763__D (.DIODE(net1564));
 sky130_fd_sc_hd__diode_2 ANTENNA__11764__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11765__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__11766__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11767__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11768__D (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11769__D (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11770__D (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11771__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11772__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11773__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11774__D (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__11775__D (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11776__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11777__D (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__11778__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__11779__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__11780__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__11781__D (.DIODE(net1444));
 sky130_fd_sc_hd__diode_2 ANTENNA__11782__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11783__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11784__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11785__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__11786__D (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11787__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__11788__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11789__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11790__D (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__CLK (.DIODE(clknet_1_1__leaf__04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11791__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11792__D (.DIODE(net1596));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__CLK (.DIODE(clknet_1_1__leaf__04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11793__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11794__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__CLK (.DIODE(clknet_1_1__leaf__04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11795__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11796__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11797__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__CLK (.DIODE(clknet_1_1__leaf__04594_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11798__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11799__D (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA__11800__D (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA__11801__D (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA__11802__D (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA__11803__D (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA__11804__D (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA__11805__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11806__D (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA__11807__D (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11808__D (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA__11809__D (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__11810__D (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA__11811__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__11812__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__11813__D (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA__11814__D (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA__11815__D (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA__11816__D (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA__11817__D (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA__11818__D (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA__11819__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__11820__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11821__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11822__D (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA__11823__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11824__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__11825__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11826__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11827__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11828__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11829__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__11830__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11831__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11832__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__11833__RESET_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__11834__RESET_B (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA__11835__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__11836__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__11837__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__11838__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__11839__D (.DIODE(net1297));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__D (.DIODE(net1574));
 sky130_fd_sc_hd__diode_2 ANTENNA__11840__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11841__D (.DIODE(net1491));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__D (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA__11842__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__D (.DIODE(net1460));
 sky130_fd_sc_hd__diode_2 ANTENNA__11843__RESET_B (.DIODE(net879));
 sky130_fd_sc_hd__diode_2 ANTENNA__11844__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__11845__D (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA__11846__D (.DIODE(net1436));
 sky130_fd_sc_hd__diode_2 ANTENNA__11847__D (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA__11848__D (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA__11849__D (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA__11850__D (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA__11851__D (.DIODE(net1508));
 sky130_fd_sc_hd__diode_2 ANTENNA__11852__D (.DIODE(net1500));
 sky130_fd_sc_hd__diode_2 ANTENNA__11853__D (.DIODE(net1484));
 sky130_fd_sc_hd__diode_2 ANTENNA__11854__D (.DIODE(net1479));
 sky130_fd_sc_hd__diode_2 ANTENNA__11855__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__11856__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__11857__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__11858__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__11859__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__11860__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__11861__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__11862__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__11863__RESET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA__11866__RESET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA__11875__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11876__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11879__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11880__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11881__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11882__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11883__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11884__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11885__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11886__CLK (.DIODE(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11887__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11888__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11889__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11890__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11891__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11892__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11893__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11894__CLK (.DIODE(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11896__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11897__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11898__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11899__RESET_B (.DIODE(net880));
 sky130_fd_sc_hd__diode_2 ANTENNA__11900__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__11901__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__11902__RESET_B (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA__11916__RESET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA__11921__RESET_B (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA__11931__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11932__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11933__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11934__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11935__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11936__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11937__CLK (.DIODE(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11938__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11939__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11940__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11941__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11942__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11943__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11944__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11945__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11946__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__11947__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11948__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11949__CLK (.DIODE(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11958__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_1[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11959__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_1[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11966__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11967__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11968__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11969__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11970__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11971__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11972__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11973__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11977__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_2[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11981__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__11982__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11983__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11984__RESET_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__11985__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11986__CLK (.DIODE(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__CLK (.DIODE(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11987__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11988__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11989__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__11990__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11991__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11992__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11993__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11994__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11995__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11996__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__CLK (.DIODE(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA__11997__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__11998__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__11999__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12000__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12001__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__12002__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__12003__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12004__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__12005__D (.DIODE(net1613));
 sky130_fd_sc_hd__diode_2 ANTENNA__12006__D (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12007__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__12008__D (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12009__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__12010__D (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12011__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12012__D (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12013__D (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA__12014__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12015__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__12016__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12017__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12018__RESET_B (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA__12019__D (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12020__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__12021__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__12022__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__12023__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__12024__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__12025__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12026__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12027__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12028__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__12029__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12030__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__12031__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12032__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12033__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__12034__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__12035__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12036__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__12037__D (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA__12038__D (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12039__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__12040__D (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12041__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__12042__D (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12043__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12044__D (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12045__D (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA__12046__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12047__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__12048__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12049__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__12050__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12051__D (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12052__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__12053__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__12054__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__12055__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__12056__D (.DIODE(net1588));
 sky130_fd_sc_hd__diode_2 ANTENNA__12057__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12058__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12059__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12060__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__12061__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12062__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__12063__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12064__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12065__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__12066__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__12067__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12068__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__12069__D (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA__12070__D (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12071__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__12072__D (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12073__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__12074__D (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12075__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12076__D (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12077__D (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA__12078__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12079__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__12080__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12081__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__12082__D (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA__12083__D (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12084__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__12085__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__12086__D (.DIODE(net1605));
 sky130_fd_sc_hd__diode_2 ANTENNA__12087__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__12088__D (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA__12089__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12090__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12091__D (.DIODE(net1558));
 sky130_fd_sc_hd__diode_2 ANTENNA__12092__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__12093__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12094__D (.DIODE(net1428));
 sky130_fd_sc_hd__diode_2 ANTENNA__12095__D (.DIODE(net1421));
 sky130_fd_sc_hd__diode_2 ANTENNA__12096__D (.DIODE(net1289));
 sky130_fd_sc_hd__diode_2 ANTENNA__12097__D (.DIODE(net1646));
 sky130_fd_sc_hd__diode_2 ANTENNA__12098__D (.DIODE(net1639));
 sky130_fd_sc_hd__diode_2 ANTENNA__12099__D (.DIODE(net1631));
 sky130_fd_sc_hd__diode_2 ANTENNA__12100__D (.DIODE(net1624));
 sky130_fd_sc_hd__diode_2 ANTENNA__12101__D (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA__12102__D (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA__12103__D (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA__12104__D (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA__12105__D (.DIODE(net1468));
 sky130_fd_sc_hd__diode_2 ANTENNA__12106__D (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA__12107__D (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA__12108__D (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA__12109__D (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA__12110__D (.DIODE(net1536));
 sky130_fd_sc_hd__diode_2 ANTENNA__12111__D (.DIODE(net1528));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__D (.DIODE(net1521));
 sky130_fd_sc_hd__diode_2 ANTENNA__12112__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12113__D (.DIODE(net1514));
 sky130_fd_sc_hd__diode_2 ANTENNA__12114__D (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA__12115__D (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA__12116__D (.DIODE(net1483));
 sky130_fd_sc_hd__diode_2 ANTENNA__12117__D (.DIODE(net1476));
 sky130_fd_sc_hd__diode_2 ANTENNA__12118__D (.DIODE(net1612));
 sky130_fd_sc_hd__diode_2 ANTENNA__12119__D (.DIODE(net1597));
 sky130_fd_sc_hd__diode_2 ANTENNA__12120__D (.DIODE(net1594));
 sky130_fd_sc_hd__diode_2 ANTENNA__12121__D (.DIODE(net1580));
 sky130_fd_sc_hd__diode_2 ANTENNA__12122__D (.DIODE(net1565));
 sky130_fd_sc_hd__diode_2 ANTENNA__12123__D (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA__12124__D (.DIODE(net1551));
 sky130_fd_sc_hd__diode_2 ANTENNA__12125__D (.DIODE(net1544));
 sky130_fd_sc_hd__diode_2 ANTENNA__12134__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12135__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12136__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12137__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12138__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12139__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12140__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12141__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12143__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12148__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12149__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12150__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12151__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12152__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12153__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12154__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12155__CLK (.DIODE(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12156__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__CLK (.DIODE(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12157__D (.DIODE(\u_pwm.u_pwm_2.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__CLK (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12158__D (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12159__RESET_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12160__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12161__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12162__RESET_B (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA__12163__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12164__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12165__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12166__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12167__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12168__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12169__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12170__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12171__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12172__RESET_B (.DIODE(net816));
 sky130_fd_sc_hd__diode_2 ANTENNA__12173__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12174__RESET_B (.DIODE(net818));
 sky130_fd_sc_hd__diode_2 ANTENNA__12176__RESET_B (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA__12181__RESET_B (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA__12231__A (.DIODE(\u_glbl_reg.reg_2[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12232__A (.DIODE(\u_glbl_reg.reg_2[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12233__A (.DIODE(\u_glbl_reg.reg_2[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12234__A (.DIODE(\u_glbl_reg.reg_2[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12235__A (.DIODE(\u_glbl_reg.reg_2[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12236__A (.DIODE(\u_glbl_reg.reg_2[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12237__A (.DIODE(\u_glbl_reg.reg_2[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12238__A (.DIODE(\u_glbl_reg.reg_2[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12239__A (.DIODE(\u_glbl_reg.reg_2[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12240__A (.DIODE(\u_glbl_reg.reg_2[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12243__A (.DIODE(\u_glbl_reg.reg_2[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12245__A (.DIODE(\u_glbl_reg.reg_2[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12246__A (.DIODE(\u_glbl_reg.reg_2[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12251__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12252__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12253__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12254__A (.DIODE(net1652));
 sky130_fd_sc_hd__diode_2 ANTENNA__12255__A (.DIODE(net1653));
 sky130_fd_sc_hd__diode_2 ANTENNA__12256__A (.DIODE(net1653));
 sky130_fd_sc_hd__diode_2 ANTENNA__12267__A (.DIODE(net1339));
 sky130_fd_sc_hd__diode_2 ANTENNA__12268__A (.DIODE(net1376));
 sky130_fd_sc_hd__diode_2 ANTENNA__12269__A (.DIODE(net1373));
 sky130_fd_sc_hd__diode_2 ANTENNA__12270__A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA__12271__A (.DIODE(net1357));
 sky130_fd_sc_hd__diode_2 ANTENNA__12272__A (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA__12273__A (.DIODE(net1345));
 sky130_fd_sc_hd__diode_2 ANTENNA__12274__A (.DIODE(net1344));
 sky130_fd_sc_hd__diode_2 ANTENNA__12275__A (.DIODE(net1342));
 sky130_fd_sc_hd__diode_2 ANTENNA__12276__A (.DIODE(net1341));
 sky130_fd_sc_hd__diode_2 ANTENNA__12277__A (.DIODE(net1340));
 sky130_fd_sc_hd__diode_2 ANTENNA__12278__A (.DIODE(net1374));
 sky130_fd_sc_hd__diode_2 ANTENNA__12279__A (.DIODE(net1337));
 sky130_fd_sc_hd__diode_2 ANTENNA__12280__A (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA__12281__A (.DIODE(net1322));
 sky130_fd_sc_hd__diode_2 ANTENNA__12282__A (.DIODE(net1315));
 sky130_fd_sc_hd__diode_2 ANTENNA__12283__A (.DIODE(net1302));
 sky130_fd_sc_hd__diode_2 ANTENNA__12284__A (.DIODE(net1576));
 sky130_fd_sc_hd__diode_2 ANTENNA__12285__A (.DIODE(net1495));
 sky130_fd_sc_hd__diode_2 ANTENNA__12286__A (.DIODE(net1472));
 sky130_fd_sc_hd__diode_2 ANTENNA__12287__A (.DIODE(net1462));
 sky130_fd_sc_hd__diode_2 ANTENNA__12288__A (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA__12289__A (.DIODE(net1446));
 sky130_fd_sc_hd__diode_2 ANTENNA__12290__A (.DIODE(net1437));
 sky130_fd_sc_hd__diode_2 ANTENNA__12291__A (.DIODE(net1431));
 sky130_fd_sc_hd__diode_2 ANTENNA__12292__A (.DIODE(net1424));
 sky130_fd_sc_hd__diode_2 ANTENNA__12293__A (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA__12294__A (.DIODE(net1649));
 sky130_fd_sc_hd__diode_2 ANTENNA__12295__A (.DIODE(net1642));
 sky130_fd_sc_hd__diode_2 ANTENNA__12296__A (.DIODE(net1634));
 sky130_fd_sc_hd__diode_2 ANTENNA__12297__A (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA__12298__A (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA__12299__A (.DIODE(net1609));
 sky130_fd_sc_hd__diode_2 ANTENNA__12300__A (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA__12301__A (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA__12302__A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA__12303__A (.DIODE(net1570));
 sky130_fd_sc_hd__diode_2 ANTENNA__12304__A (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA__12305__A (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA__12306__A (.DIODE(net1548));
 sky130_fd_sc_hd__diode_2 ANTENNA__12307__A (.DIODE(net1540));
 sky130_fd_sc_hd__diode_2 ANTENNA__12308__A (.DIODE(net1532));
 sky130_fd_sc_hd__diode_2 ANTENNA__12309__A (.DIODE(net1525));
 sky130_fd_sc_hd__diode_2 ANTENNA__12310__A (.DIODE(net1518));
 sky130_fd_sc_hd__diode_2 ANTENNA__12311__A (.DIODE(net1511));
 sky130_fd_sc_hd__diode_2 ANTENNA__12312__A (.DIODE(net1504));
 sky130_fd_sc_hd__diode_2 ANTENNA__12313__A (.DIODE(net1487));
 sky130_fd_sc_hd__diode_2 ANTENNA__12314__A (.DIODE(net1480));
 sky130_fd_sc_hd__diode_2 ANTENNA__12315__A (.DIODE(net1416));
 sky130_fd_sc_hd__diode_2 ANTENNA__12316__A (.DIODE(net1395));
 sky130_fd_sc_hd__diode_2 ANTENNA__12317__A (.DIODE(net1393));
 sky130_fd_sc_hd__diode_2 ANTENNA__12318__A (.DIODE(net1391));
 sky130_fd_sc_hd__diode_2 ANTENNA__12319__A (.DIODE(net1389));
 sky130_fd_sc_hd__diode_2 ANTENNA__12320__A (.DIODE(\u_glbl_reg.reg_12[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12324__A (.DIODE(\u_glbl_reg.reg_2[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12326__A (.DIODE(\u_glbl_reg.reg_2[2] ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12327__A (.DIODE(net1375));
 sky130_fd_sc_hd__diode_2 ANTENNA__12333__GATE (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12334__GATE (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12375__CLK (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12381__CLK (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12414__CLK (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12421__CLK (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12440__GATE (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12441__GATE (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA__12442__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12443__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12444__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12445__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12446__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12447__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12448__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12449__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12450__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12451__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12452__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12453__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12454__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12455__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12456__GATE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__12457__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12458__GATE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__12459__GATE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__12460__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12461__GATE (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12462__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12463__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12464__GATE (.DIODE(net719));
 sky130_fd_sc_hd__diode_2 ANTENNA__12465__GATE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__12466__GATE (.DIODE(net722));
 sky130_fd_sc_hd__diode_2 ANTENNA__12467__GATE (.DIODE(net721));
 sky130_fd_sc_hd__diode_2 ANTENNA__12488__CLK (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12523__CLK (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12531__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12532__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12533__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12534__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12535__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12536__GATE (.DIODE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12547__CLK (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12555__CLK (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12557__CLK (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12559__GATE (.DIODE(_00403_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12573__CLK (.DIODE(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12583__GATE (.DIODE(_00458_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12584__GATE (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12585__GATE (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12586__GATE (.DIODE(_00459_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12601__CLK (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12606__GATE (.DIODE(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__diode_2 ANTENNA__12607__GATE (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA__12615__CLK (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12620__CLK (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12635__GATE (.DIODE(_00589_));
 sky130_fd_sc_hd__diode_2 ANTENNA__12645__CLK (.DIODE(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12648__CLK (.DIODE(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA__12654__CLK (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04353__A (.DIODE(_04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04358__A (.DIODE(_04358_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04359__A (.DIODE(_04359_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04406__A (.DIODE(_04406_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04493__A (.DIODE(_04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04586__A (.DIODE(_04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04587__A (.DIODE(_04587_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04589__A (.DIODE(_04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0__04608__A (.DIODE(_04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_mclk_A (.DIODE(net1692));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock1_A (.DIODE(user_clock1));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_0_user_clock2_A (.DIODE(user_clock2));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0_0_mclk_A (.DIODE(net1695));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04353__A (.DIODE(clknet_0__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04493__A (.DIODE(clknet_0__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04564__A (.DIODE(clknet_0__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04567__A (.DIODE(clknet_0__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04586__A (.DIODE(clknet_0__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04589__A (.DIODE(clknet_0__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04608__A (.DIODE(clknet_0__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_0__f__04611__A (.DIODE(clknet_0__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1_0_mclk_A (.DIODE(clknet_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04353__A (.DIODE(clknet_0__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04493__A (.DIODE(clknet_0__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04564__A (.DIODE(clknet_0__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04567__A (.DIODE(clknet_0__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04586__A (.DIODE(clknet_0__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04589__A (.DIODE(clknet_0__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04608__A (.DIODE(clknet_0__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_1__f__04611__A (.DIODE(clknet_0__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2_0_mclk_A (.DIODE(net1696));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04353__A (.DIODE(clknet_0__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04493__A (.DIODE(clknet_0__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04564__A (.DIODE(clknet_0__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04567__A (.DIODE(clknet_0__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04586__A (.DIODE(clknet_0__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04589__A (.DIODE(clknet_0__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04608__A (.DIODE(clknet_0__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_2__f__04611__A (.DIODE(clknet_0__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3_0_mclk_A (.DIODE(net1696));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04353__A (.DIODE(clknet_0__04353_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04493__A (.DIODE(clknet_0__04493_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04564__A (.DIODE(clknet_0__04564_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04567__A (.DIODE(clknet_0__04567_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04586__A (.DIODE(clknet_0__04586_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04589__A (.DIODE(clknet_0__04589_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04608__A (.DIODE(clknet_0__04608_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_2_3__f__04611__A (.DIODE(clknet_0__04611_));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_0__f_mclk_A (.DIODE(clknet_2_0_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_10__f_mclk_A (.DIODE(clknet_2_2_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_11__f_mclk_A (.DIODE(clknet_2_2_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_12__f_mclk_A (.DIODE(clknet_2_3_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_13__f_mclk_A (.DIODE(clknet_2_3_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_14__f_mclk_A (.DIODE(clknet_2_3_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_15__f_mclk_A (.DIODE(clknet_2_3_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_1__f_mclk_A (.DIODE(clknet_2_0_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_2__f_mclk_A (.DIODE(clknet_2_0_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_3__f_mclk_A (.DIODE(clknet_2_0_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_4__f_mclk_A (.DIODE(clknet_2_1_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_5__f_mclk_A (.DIODE(clknet_2_1_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_6__f_mclk_A (.DIODE(clknet_2_1_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_7__f_mclk_A (.DIODE(clknet_2_1_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_8__f_mclk_A (.DIODE(clknet_2_2_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_4_9__f_mclk_A (.DIODE(clknet_2_2_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_0_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_100_mclk_A (.DIODE(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_102_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_103_mclk_A (.DIODE(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_104_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_105_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_106_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_107_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_109_mclk_A (.DIODE(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_10_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_110_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_111_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_112_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_113_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_114_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_115_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_116_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_117_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_118_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_11_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_120_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_122_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_123_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_124_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_126_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_127_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_128_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_12_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_13_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_14_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_15_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_16_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_17_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_19_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_1_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_20_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_21_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_22_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_23_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_24_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_25_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_26_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_28_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_29_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_2_mclk_A (.DIODE(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_30_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_31_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_32_mclk_A (.DIODE(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_33_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_34_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_35_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_36_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_37_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_38_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_39_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_40_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_41_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_42_mclk_A (.DIODE(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_43_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_44_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_45_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_46_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_47_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_48_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_4_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_51_mclk_A (.DIODE(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_53_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_54_mclk_A (.DIODE(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_55_mclk_A (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_56_mclk_A (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_58_mclk_A (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_5_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_60_mclk_A (.DIODE(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_62_mclk_A (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_63_mclk_A (.DIODE(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_65_mclk_A (.DIODE(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_66_mclk_A (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_67_mclk_A (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_69_mclk_A (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_6_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_70_mclk_A (.DIODE(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_72_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_73_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_74_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_75_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_76_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_77_mclk_A (.DIODE(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_78_mclk_A (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_79_mclk_A (.DIODE(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_7_mclk_A (.DIODE(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_80_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_81_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_82_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_83_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_84_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_85_mclk_A (.DIODE(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_86_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_87_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_88_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_89_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_8_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_90_mclk_A (.DIODE(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_91_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_92_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_93_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_94_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_95_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_96_mclk_A (.DIODE(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_97_mclk_A (.DIODE(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_99_mclk_A (.DIODE(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_clkbuf_leaf_9_mclk_A (.DIODE(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1002_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1006_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1007_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1010_A (.DIODE(net1011));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1011_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1013_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1015_A (.DIODE(net1016));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1016_A (.DIODE(net1017));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1017_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1018_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1020_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1021_A (.DIODE(net1022));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1022_A (.DIODE(net1023));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1023_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1025_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1026_A (.DIODE(net1027));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1027_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1028_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1029_A (.DIODE(net1030));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1030_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1031_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1032_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1034_A (.DIODE(net1035));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1035_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1036_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1037_A (.DIODE(net1038));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1039_A (.DIODE(net1040));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1040_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1041_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1044_A (.DIODE(net1045));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1045_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1046_A (.DIODE(net1047));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1047_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1048_A (.DIODE(net1049));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1049_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1050_A (.DIODE(net1051));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1051_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1052_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1053_A (.DIODE(net1054));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1054_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1055_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1056_A (.DIODE(net1057));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1057_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1058_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1059_A (.DIODE(net1060));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1060_A (.DIODE(net1061));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1062_A (.DIODE(net1063));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1063_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1064_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1065_A (.DIODE(net1066));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1067_A (.DIODE(net1069));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1074_A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1075_A (.DIODE(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1080_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1081_A (.DIODE(net1082));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1083_A (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1084_A (.DIODE(net1085));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1086_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1087_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1088_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1089_A (.DIODE(net1090));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1091_A (.DIODE(\reg_blk_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1092_A (.DIODE(\reg_blk_sel[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1109_A (.DIODE(\u_glbl_reg.cfg_multi_func_sel[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1110_A (.DIODE(_03462_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1111_A (.DIODE(net1112));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1112_A (.DIODE(net1113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1114_A (.DIODE(net1115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1115_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1116_A (.DIODE(net1117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1117_A (.DIODE(net1118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1119_A (.DIODE(net1120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1120_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1121_A (.DIODE(net1122));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1122_A (.DIODE(net1123));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1124_A (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1125_A (.DIODE(net1126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1126_A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1127_A (.DIODE(net1128));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1128_A (.DIODE(_01546_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1131_A (.DIODE(net1132));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1132_A (.DIODE(net1133));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1133_A (.DIODE(_01541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1134_A (.DIODE(_01541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1135_A (.DIODE(_01541_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1136_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1137_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1138_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1139_A (.DIODE(net1140));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1140_A (.DIODE(net1141));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1142_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1143_A (.DIODE(net1144));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1144_A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1145_A (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1146_A (.DIODE(net1147));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1147_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1149_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1150_A (.DIODE(net1151));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1151_A (.DIODE(_01349_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1152_A (.DIODE(net1153));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1154_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1155_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1156_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1157_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1158_A (.DIODE(net1159));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1159_A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1160_A (.DIODE(net1161));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1161_A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1162_A (.DIODE(net1163));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1163_A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1164_A (.DIODE(net1165));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1165_A (.DIODE(_01114_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1166_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1167_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1168_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1169_A (.DIODE(net1170));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1170_A (.DIODE(net1171));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1171_A (.DIODE(_01113_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1172_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1173_A (.DIODE(net1174));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1174_A (.DIODE(_01113_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1175_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1176_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1177_A (.DIODE(net1178));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1179_A (.DIODE(_00998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1180_A (.DIODE(_00998_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1181_A (.DIODE(net1182));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1182_A (.DIODE(_00996_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1201_A (.DIODE(net1202));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1202_A (.DIODE(net2293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1203_A (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1204_A (.DIODE(net1205));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1205_A (.DIODE(net2293));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1207_A (.DIODE(net1208));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1208_A (.DIODE(net1209));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1209_A (.DIODE(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1210_A (.DIODE(net1729));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1211_A (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1212_A (.DIODE(net1213));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1214_A (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1215_A (.DIODE(net1216));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1216_A (.DIODE(_01129_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1217_A (.DIODE(net1218));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1218_A (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1219_A (.DIODE(net1220));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1220_A (.DIODE(net1221));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1221_A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1222_A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1223_A (.DIODE(net1224));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1224_A (.DIODE(net1225));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1226_A (.DIODE(net1227));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1227_A (.DIODE(net1228));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1228_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1229_A (.DIODE(net1230));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1230_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1231_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1232_A (.DIODE(net1233));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1234_A (.DIODE(net1235));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1235_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1236_A (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1237_A (.DIODE(net1238));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1238_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1239_A (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1240_A (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1241_A (.DIODE(net1242));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1242_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1243_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1244_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1245_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1246_A (.DIODE(net1247));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1247_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1248_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1249_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1250_A (.DIODE(net1251));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1251_A (.DIODE(net1252));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1252_A (.DIODE(net1253));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1254_A (.DIODE(net1255));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1256_A (.DIODE(net1257));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1257_A (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1258_A (.DIODE(net1259));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1259_A (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1260_A (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1261_A (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1262_A (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1263_A (.DIODE(net1264));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1264_A (.DIODE(net1265));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1266_A (.DIODE(net1267));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1267_A (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1268_A (.DIODE(net1269));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1269_A (.DIODE(net1270));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1270_A (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1271_A (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1272_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1273_A (.DIODE(net1274));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1274_A (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1275_A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1276_A (.DIODE(net1277));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1277_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1278_A (.DIODE(net1279));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1279_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1280_A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1281_A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1282_A (.DIODE(net1283));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1283_A (.DIODE(net1285));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1286_A (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1287_A (.DIODE(net1288));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1288_A (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1289_A (.DIODE(net1290));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1291_A (.DIODE(net1292));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1293_A (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1294_A (.DIODE(net1295));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1295_A (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1296_A (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1297_A (.DIODE(net1298));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1298_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1299_A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1300_A (.DIODE(net1301));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1301_A (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1302_A (.DIODE(net1303));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1303_A (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1308_A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1309_A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1310_A (.DIODE(net1311));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1312_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1316_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1317_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1319_A (.DIODE(net1320));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1320_A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1321_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1323_A (.DIODE(net1325));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1324_A (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1325_A (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1326_A (.DIODE(net1328));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1329_A (.DIODE(net1330));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1331_A (.DIODE(net1332));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1332_A (.DIODE(net1333));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1333_A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1334_A (.DIODE(net1335));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1335_A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1336_A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1337_A (.DIODE(net1338));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1343_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1344_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1346_A (.DIODE(net1347));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1348_A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1349_A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1350_A (.DIODE(net1351));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1351_A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1352_A (.DIODE(net1353));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1353_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1354_A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1355_A (.DIODE(net1356));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1356_A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1357_A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1358_A (.DIODE(net1359));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1359_A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1360_A (.DIODE(net1361));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1361_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1362_A (.DIODE(net1363));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1363_A (.DIODE(net1364));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1364_A (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1366_A (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1367_A (.DIODE(net1368));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1368_A (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1369_A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1370_A (.DIODE(net1371));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1371_A (.DIODE(net1372));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1372_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1378_A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1379_A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1380_A (.DIODE(net1381));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1381_A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1382_A (.DIODE(net1383));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1383_A (.DIODE(net1384));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1384_A (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1385_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1418_A (.DIODE(net1419));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1419_A (.DIODE(net1420));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1420_A (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1421_A (.DIODE(net1422));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1423_A (.DIODE(net1424));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1425_A (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1426_A (.DIODE(net1427));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1428_A (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1429_A (.DIODE(net1431));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1433_A (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1434_A (.DIODE(net1435));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1435_A (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1436_A (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1437_A (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1438_A (.DIODE(net1440));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1440_A (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1441_A (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1442_A (.DIODE(net1443));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1443_A (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1444_A (.DIODE(net1445));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1445_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1446_A (.DIODE(net1447));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1447_A (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1448_A (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1449_A (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1450_A (.DIODE(net1451));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1451_A (.DIODE(net1452));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1452_A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1453_A (.DIODE(net1455));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1454_A (.DIODE(net1456));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1457_A (.DIODE(net1458));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1458_A (.DIODE(net1459));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1459_A (.DIODE(net1465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1460_A (.DIODE(net1461));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1461_A (.DIODE(net1465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1463_A (.DIODE(net1465));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1466_A (.DIODE(net1467));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1467_A (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1468_A (.DIODE(net1469));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1469_A (.DIODE(net1473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1471_A (.DIODE(net1473));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1474_A (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1475_A (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1476_A (.DIODE(net1477));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1477_A (.DIODE(net1478));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1478_A (.DIODE(net1479));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1481_A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1482_A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1483_A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1484_A (.DIODE(net1485));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1485_A (.DIODE(net1486));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1486_A (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1488_A (.DIODE(net1489));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1489_A (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1490_A (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1491_A (.DIODE(net1492));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1492_A (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1493_A (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1494_A (.DIODE(net1496));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1496_A (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1498_A (.DIODE(net1499));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1499_A (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1500_A (.DIODE(net1501));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1501_A (.DIODE(net1502));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1503_A (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1505_A (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1506_A (.DIODE(net1507));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1507_A (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1508_A (.DIODE(net1509));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1509_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1510_A (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1512_A (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1513_A (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1514_A (.DIODE(net1515));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1515_A (.DIODE(net1516));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1516_A (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1517_A (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1519_A (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1520_A (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1521_A (.DIODE(net1522));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1522_A (.DIODE(net1523));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1523_A (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1526_A (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1527_A (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1528_A (.DIODE(net1529));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1529_A (.DIODE(net1530));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1531_A (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1534_A (.DIODE(net1535));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1535_A (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1536_A (.DIODE(net1537));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1537_A (.DIODE(net1538));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1538_A (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1539_A (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1541_A (.DIODE(net1542));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1543_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1545_A (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1546_A (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1547_A (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1549_A (.DIODE(net1550));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1550_A (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1551_A (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1552_A (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1553_A (.DIODE(net1554));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1554_A (.DIODE(net1555));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1556_A (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1557_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1559_A (.DIODE(net1560));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1561_A (.DIODE(net1563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1562_A (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1564_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1565_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1566_A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1567_A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1568_A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1569_A (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1572_A (.DIODE(net1573));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1573_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1574_A (.DIODE(net1575));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1575_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1576_A (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1577_A (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1579_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1580_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1581_A (.DIODE(net1582));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1583_A (.DIODE(net1585));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1584_A (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1586_A (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1587_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1589_A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1590_A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1591_A (.DIODE(net1593));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1592_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1595_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1597_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1598_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1599_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1600_A (.DIODE(net1601));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1601_A (.DIODE(net1602));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1603_A (.DIODE(net1604));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1606_A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1608_A (.DIODE(net1611));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1613_A (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1614_A (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1615_A (.DIODE(net1616));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1616_A (.DIODE(net1617));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1618_A (.DIODE(net1620));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1621_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1622_A (.DIODE(net1623));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1623_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1624_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1625_A (.DIODE(net1627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1628_A (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1629_A (.DIODE(net1630));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1631_A (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1632_A (.DIODE(net1634));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1636_A (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1637_A (.DIODE(net1638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1638_A (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1639_A (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1640_A (.DIODE(net1642));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1643_A (.DIODE(net1644));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1644_A (.DIODE(net1645));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1645_A (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1646_A (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1647_A (.DIODE(net1649));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout1651_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout517_A (.DIODE(net518));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout518_A (.DIODE(_04039_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout519_A (.DIODE(_01348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout520_A (.DIODE(_01348_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout521_A (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout522_A (.DIODE(_01343_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout541_A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout542_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout543_A (.DIODE(net544));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout544_A (.DIODE(net545));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout546_A (.DIODE(net547));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout547_A (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout548_A (.DIODE(_03475_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout549_A (.DIODE(_03472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout550_A (.DIODE(_03472_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout552_A (.DIODE(_03471_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout553_A (.DIODE(_03470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout554_A (.DIODE(_03470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout555_A (.DIODE(_03470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout556_A (.DIODE(_03470_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout557_A (.DIODE(net558));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout559_A (.DIODE(_03464_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout560_A (.DIODE(net561));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout561_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout562_A (.DIODE(net563));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout563_A (.DIODE(_01785_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout573_A (.DIODE(net574));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout574_A (.DIODE(_01198_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout575_A (.DIODE(_01005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout576_A (.DIODE(_01005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout577_A (.DIODE(net578));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout578_A (.DIODE(_01005_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout584_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout585_A (.DIODE(net586));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout589_A (.DIODE(net590));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout590_A (.DIODE(_01793_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout591_A (.DIODE(_01793_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout592_A (.DIODE(_01793_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout593_A (.DIODE(net594));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout594_A (.DIODE(net595));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout596_A (.DIODE(_01782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout597_A (.DIODE(_01782_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout598_A (.DIODE(net599));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout599_A (.DIODE(net600));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout603_A (.DIODE(net604));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout604_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout605_A (.DIODE(net606));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout607_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout608_A (.DIODE(net609));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout609_A (.DIODE(_01557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout610_A (.DIODE(_01557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout611_A (.DIODE(_01557_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout612_A (.DIODE(net613));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout613_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout614_A (.DIODE(net615));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout616_A (.DIODE(net617));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout617_A (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout618_A (.DIODE(net619));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout620_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout621_A (.DIODE(net622));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout622_A (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout623_A (.DIODE(_01554_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout624_A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout625_A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout626_A (.DIODE(net627));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout627_A (.DIODE(_01553_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout628_A (.DIODE(net629));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout629_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout630_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout631_A (.DIODE(net632));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout632_A (.DIODE(_01552_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout633_A (.DIODE(net634));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout634_A (.DIODE(_01551_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout635_A (.DIODE(net636));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout636_A (.DIODE(_01551_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout637_A (.DIODE(net638));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout638_A (.DIODE(_01550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout639_A (.DIODE(_01550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout640_A (.DIODE(_01550_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout641_A (.DIODE(net642));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout642_A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout643_A (.DIODE(net644));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout645_A (.DIODE(_01548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout646_A (.DIODE(_01548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout647_A (.DIODE(net648));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout648_A (.DIODE(_01548_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout649_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout650_A (.DIODE(net651));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout651_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout652_A (.DIODE(net653));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout653_A (.DIODE(_01547_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout654_A (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout655_A (.DIODE(net656));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout656_A (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout657_A (.DIODE(net658));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout658_A (.DIODE(_01545_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout659_A (.DIODE(net660));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout660_A (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout661_A (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout662_A (.DIODE(net663));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout664_A (.DIODE(net665));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout665_A (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout666_A (.DIODE(net667));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout667_A (.DIODE(_01539_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout668_A (.DIODE(net669));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout669_A (.DIODE(_01538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout670_A (.DIODE(_01538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout671_A (.DIODE(_01538_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout672_A (.DIODE(net673));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout674_A (.DIODE(_01482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout675_A (.DIODE(_01482_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout676_A (.DIODE(_01463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout677_A (.DIODE(_01463_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout678_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout679_A (.DIODE(net680));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout681_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout682_A (.DIODE(net683));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout683_A (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout684_A (.DIODE(_01146_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout685_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout686_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout687_A (.DIODE(net688));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout688_A (.DIODE(net689));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout689_A (.DIODE(net690));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout690_A (.DIODE(_01134_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout691_A (.DIODE(net692));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout692_A (.DIODE(net693));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout693_A (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout694_A (.DIODE(net695));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout695_A (.DIODE(net696));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout696_A (.DIODE(net697));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout697_A (.DIODE(_01133_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout698_A (.DIODE(_01132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout699_A (.DIODE(_01132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout700_A (.DIODE(_01132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout701_A (.DIODE(_01132_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout702_A (.DIODE(net703));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout703_A (.DIODE(net704));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout704_A (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout705_A (.DIODE(net706));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout706_A (.DIODE(net707));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout707_A (.DIODE(_01131_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout708_A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout709_A (.DIODE(net710));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout710_A (.DIODE(net711));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout712_A (.DIODE(net713));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout713_A (.DIODE(net714));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout714_A (.DIODE(_01001_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout715_A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout716_A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout717_A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout718_A (.DIODE(_01000_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout719_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout720_A (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout722_A (.DIODE(_00250_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout726_A (.DIODE(_00888_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout727_A (.DIODE(_00878_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout730_A (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout731_A (.DIODE(_00837_));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout732_A (.DIODE(net733));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout733_A (.DIODE(net734));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout738_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout741_A (.DIODE(net742));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout743_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout744_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout745_A (.DIODE(net746));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout746_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout748_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout749_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout750_A (.DIODE(net751));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout751_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout755_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout758_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout762_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout763_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout764_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout765_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout766_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout767_A (.DIODE(net768));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout768_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout770_A (.DIODE(net771));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout771_A (.DIODE(net772));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout772_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout773_A (.DIODE(net774));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout774_A (.DIODE(net775));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout775_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout779_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout780_A (.DIODE(net781));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout781_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout782_A (.DIODE(net783));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout783_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout786_A (.DIODE(net787));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout788_A (.DIODE(net789));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout789_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout791_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout792_A (.DIODE(net793));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout793_A (.DIODE(net794));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout794_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout797_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout800_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout803_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout804_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout805_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout806_A (.DIODE(net807));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout807_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout808_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout809_A (.DIODE(net810));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout810_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout811_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout812_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout813_A (.DIODE(net814));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout814_A (.DIODE(net815));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout815_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout816_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout817_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout818_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout819_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout820_A (.DIODE(net821));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout821_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout825_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout826_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout828_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout829_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout830_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout831_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout834_A (.DIODE(net835));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout835_A (.DIODE(net836));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout836_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout838_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout842_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout846_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout847_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout848_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout849_A (.DIODE(net850));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout850_A (.DIODE(net851));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout851_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout855_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout856_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout857_A (.DIODE(net858));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout858_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout859_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout860_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout861_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout862_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout865_A (.DIODE(net866));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout866_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout868_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout870_A (.DIODE(net871));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout871_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout872_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout873_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout874_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout877_A (.DIODE(net878));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout878_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout879_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout880_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout881_A (.DIODE(net882));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout882_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout886_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout889_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout892_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout893_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout894_A (.DIODE(net895));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout895_A (.DIODE(net896));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout896_A (.DIODE(net897));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout897_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout898_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout899_A (.DIODE(net900));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout900_A (.DIODE(net901));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout901_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout902_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout903_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout904_A (.DIODE(net905));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout905_A (.DIODE(net906));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout906_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout907_A (.DIODE(net908));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout908_A (.DIODE(net909));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout909_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout910_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout911_A (.DIODE(net912));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout912_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout913_A (.DIODE(net914));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout914_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout915_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout916_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout917_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout918_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout919_A (.DIODE(net920));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout920_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout922_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout923_A (.DIODE(net924));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout924_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout925_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout926_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout928_A (.DIODE(net929));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout929_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout932_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout934_A (.DIODE(net935));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout935_A (.DIODE(net936));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout936_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout938_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout941_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout942_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout943_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout944_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout945_A (.DIODE(net946));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout946_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout950_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout953_A (.DIODE(net954));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout954_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout957_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout958_A (.DIODE(net959));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout959_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout964_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout967_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout968_A (.DIODE(net969));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout969_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout972_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout974_A (.DIODE(net975));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout975_A (.DIODE(net1043));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout977_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout980_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout984_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout987_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout989_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout992_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout994_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout997_A (.DIODE(net998));
 sky130_fd_sc_hd__diode_2 ANTENNA_fanout998_A (.DIODE(net1041));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold100_A (.DIODE(net436));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold103_A (.DIODE(net433));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold106_A (.DIODE(net431));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold109_A (.DIODE(_03664_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold10_A (.DIODE(net426));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold110_A (.DIODE(net437));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold113_A (.DIODE(net430));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold127_A (.DIODE(\u_pwm.u_pwm_2.cfg_pwm_run ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold153_A (.DIODE(\u_gpio.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold159_A (.DIODE(\u_glbl_reg.u_random.n1[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold165_A (.DIODE(\u_glbl_reg.u_random.n1[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold16_A (.DIODE(net427));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold172_A (.DIODE(\u_glbl_reg.u_random.n1[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold177_A (.DIODE(\u_glbl_reg.u_random.n1[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold178_A (.DIODE(\u_glbl_reg.u_random.n1[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold182_A (.DIODE(\u_glbl_reg.u_random.n0[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold183_A (.DIODE(\u_glbl_reg.u_random.n1[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold185_A (.DIODE(\u_glbl_reg.u_random.n0[17] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold186_A (.DIODE(\u_glbl_reg.u_random.n1[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold187_A (.DIODE(\u_glbl_reg.u_random.n1[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold188_A (.DIODE(\u_glbl_reg.u_random.n1[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold189_A (.DIODE(\u_glbl_reg.u_random.n1[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold190_A (.DIODE(\u_glbl_reg.u_random.n0[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold191_A (.DIODE(\u_glbl_reg.u_random.n1[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold192_A (.DIODE(\u_glbl_reg.u_random.n1[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold193_A (.DIODE(\u_glbl_reg.u_random.n0[24] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold199_A (.DIODE(\u_glbl_reg.u_random.n1[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold202_A (.DIODE(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold203_A (.DIODE(\u_glbl_reg.u_random.n1[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold204_A (.DIODE(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold205_A (.DIODE(\u_glbl_reg.u_random.n1[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold206_A (.DIODE(\u_glbl_reg.u_random.n0[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold207_A (.DIODE(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold208_A (.DIODE(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold209_A (.DIODE(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold210_A (.DIODE(\u_glbl_reg.u_random.n0[14] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold213_A (.DIODE(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold214_A (.DIODE(\u_glbl_reg.u_random.n0[31] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold215_A (.DIODE(\u_glbl_reg.u_random.n1[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold216_A (.DIODE(\u_glbl_reg.u_random.n0[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold217_A (.DIODE(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold218_A (.DIODE(\u_glbl_reg.u_random.n0[16] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold219_A (.DIODE(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold220_A (.DIODE(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold223_A (.DIODE(\u_gpio.u_bit[25].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold227_A (.DIODE(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold228_A (.DIODE(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold229_A (.DIODE(\u_glbl_reg.u_random.n0[22] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold230_A (.DIODE(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold231_A (.DIODE(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold232_A (.DIODE(\u_glbl_reg.u_random.n0[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold233_A (.DIODE(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold240_A (.DIODE(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold241_A (.DIODE(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold266_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold268_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold283_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold28_A (.DIODE(net425));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold291_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold302_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold30_A (.DIODE(\u_pwm.blk_sel[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold314_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold315_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold326_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold336_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold357_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold364_A (.DIODE(\u_glbl_reg.reg_out[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold366_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold367_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold392_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold395_A (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold398_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold3_A (.DIODE(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold427_A (.DIODE(\u_pwm.u_pwm_0.u_reg.reg_2[18] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold43_A (.DIODE(net429));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold46_A (.DIODE(net418));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold49_A (.DIODE(net440));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold524_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold52_A (.DIODE(net443));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold548_A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold55_A (.DIODE(net444));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold58_A (.DIODE(net445));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold603_A (.DIODE(\u_ws281x.u_reg.gfifo[1].u_fifo.full ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold618_A (.DIODE(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold619_A (.DIODE(\u_glbl_reg.reg_out[0] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold61_A (.DIODE(net449));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold630_A (.DIODE(\u_ws281x.port1_enb ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold64_A (.DIODE(net419));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold67_A (.DIODE(net442));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(\u_glbl_reg.cfg_rst_ctrl[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold70_A (.DIODE(net448));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold75_A (.DIODE(net441));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold78_A (.DIODE(_03676_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold79_A (.DIODE(net439));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold82_A (.DIODE(_03652_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold83_A (.DIODE(net435));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold86_A (.DIODE(_03634_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold87_A (.DIODE(net432));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold90_A (.DIODE(net434));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold92_A (.DIODE(\u_glbl_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold93_A (.DIODE(net438));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold96_A (.DIODE(_03616_));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold97_A (.DIODE(net428));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold99_A (.DIODE(\u_glbl_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_input100_A (.DIODE(reg_wdata[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input101_A (.DIODE(reg_wdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input102_A (.DIODE(reg_wdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input103_A (.DIODE(reg_wdata[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input104_A (.DIODE(reg_wdata[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input105_A (.DIODE(reg_wdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input106_A (.DIODE(reg_wdata[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input107_A (.DIODE(reg_wdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input108_A (.DIODE(reg_wdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input109_A (.DIODE(reg_wdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input10_A (.DIODE(digital_io_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input110_A (.DIODE(reg_wdata[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input111_A (.DIODE(reg_wdata[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input112_A (.DIODE(reg_wdata[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input113_A (.DIODE(reg_wdata[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input114_A (.DIODE(reg_wdata[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input115_A (.DIODE(reg_wdata[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input116_A (.DIODE(reg_wdata[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input117_A (.DIODE(reg_wdata[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input118_A (.DIODE(reg_wdata[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input119_A (.DIODE(reg_wdata[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input11_A (.DIODE(digital_io_in[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input120_A (.DIODE(reg_wdata[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input121_A (.DIODE(reg_wdata[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input122_A (.DIODE(reg_wdata[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input123_A (.DIODE(reg_wdata[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input124_A (.DIODE(reg_wdata[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input125_A (.DIODE(reg_wdata[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input126_A (.DIODE(reg_wdata[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input127_A (.DIODE(reg_wdata[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input128_A (.DIODE(reg_wdata[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input129_A (.DIODE(reg_wdata[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input12_A (.DIODE(digital_io_in[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input130_A (.DIODE(reg_wr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input131_A (.DIODE(riscv_tdo));
 sky130_fd_sc_hd__diode_2 ANTENNA_input132_A (.DIODE(riscv_tdo_en));
 sky130_fd_sc_hd__diode_2 ANTENNA_input133_A (.DIODE(rtc_intr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input134_A (.DIODE(s_reset_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input135_A (.DIODE(sflash_do[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input136_A (.DIODE(sflash_do[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input137_A (.DIODE(sflash_do[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input138_A (.DIODE(sflash_do[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input139_A (.DIODE(sflash_oen[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input13_A (.DIODE(digital_io_in[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input140_A (.DIODE(sflash_oen[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input141_A (.DIODE(sflash_oen[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input142_A (.DIODE(sflash_oen[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input143_A (.DIODE(sflash_sck));
 sky130_fd_sc_hd__diode_2 ANTENNA_input144_A (.DIODE(sflash_ss[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input145_A (.DIODE(sflash_ss[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input146_A (.DIODE(sflash_ss[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input147_A (.DIODE(sflash_ss[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input148_A (.DIODE(sm_a1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input149_A (.DIODE(sm_a2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input14_A (.DIODE(digital_io_in[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input150_A (.DIODE(sm_b1));
 sky130_fd_sc_hd__diode_2 ANTENNA_input151_A (.DIODE(sm_b2));
 sky130_fd_sc_hd__diode_2 ANTENNA_input152_A (.DIODE(spim_miso));
 sky130_fd_sc_hd__diode_2 ANTENNA_input153_A (.DIODE(spim_sck));
 sky130_fd_sc_hd__diode_2 ANTENNA_input154_A (.DIODE(spim_ssn[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input155_A (.DIODE(spim_ssn[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input156_A (.DIODE(spim_ssn[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input157_A (.DIODE(spim_ssn[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input158_A (.DIODE(spis_miso));
 sky130_fd_sc_hd__diode_2 ANTENNA_input159_A (.DIODE(system_strap[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input15_A (.DIODE(digital_io_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input160_A (.DIODE(system_strap[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input161_A (.DIODE(system_strap[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input162_A (.DIODE(system_strap[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input163_A (.DIODE(system_strap[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input164_A (.DIODE(system_strap[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input165_A (.DIODE(system_strap[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input166_A (.DIODE(system_strap[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input167_A (.DIODE(system_strap[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input168_A (.DIODE(system_strap[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input169_A (.DIODE(system_strap[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input16_A (.DIODE(digital_io_in[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input170_A (.DIODE(system_strap[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input171_A (.DIODE(system_strap[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input172_A (.DIODE(system_strap[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input173_A (.DIODE(system_strap[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input174_A (.DIODE(system_strap[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input175_A (.DIODE(system_strap[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input176_A (.DIODE(system_strap[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input177_A (.DIODE(system_strap[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input178_A (.DIODE(system_strap[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input179_A (.DIODE(system_strap[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input17_A (.DIODE(digital_io_in[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input180_A (.DIODE(system_strap[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input181_A (.DIODE(system_strap[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input182_A (.DIODE(system_strap[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input183_A (.DIODE(system_strap[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input184_A (.DIODE(system_strap[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input185_A (.DIODE(system_strap[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input186_A (.DIODE(system_strap[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input187_A (.DIODE(system_strap[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input188_A (.DIODE(system_strap[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input189_A (.DIODE(system_strap[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input18_A (.DIODE(digital_io_in[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input190_A (.DIODE(system_strap[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input191_A (.DIODE(uart_txd[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input192_A (.DIODE(uart_txd[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input193_A (.DIODE(uartm_txd));
 sky130_fd_sc_hd__diode_2 ANTENNA_input194_A (.DIODE(usb_dn_o));
 sky130_fd_sc_hd__diode_2 ANTENNA_input195_A (.DIODE(usb_dp_o));
 sky130_fd_sc_hd__diode_2 ANTENNA_input196_A (.DIODE(usb_intr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input197_A (.DIODE(usb_oen));
 sky130_fd_sc_hd__diode_2 ANTENNA_input198_A (.DIODE(wbd_clk_int));
 sky130_fd_sc_hd__diode_2 ANTENNA_input19_A (.DIODE(digital_io_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input1_A (.DIODE(cfg_strap_pad_ctrl));
 sky130_fd_sc_hd__diode_2 ANTENNA_input20_A (.DIODE(digital_io_in[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input21_A (.DIODE(digital_io_in[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input22_A (.DIODE(digital_io_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input23_A (.DIODE(digital_io_in[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input24_A (.DIODE(digital_io_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input25_A (.DIODE(digital_io_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input26_A (.DIODE(digital_io_in[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input27_A (.DIODE(digital_io_in[32]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input28_A (.DIODE(digital_io_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input29_A (.DIODE(digital_io_in[34]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input2_A (.DIODE(cpu_clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_input30_A (.DIODE(digital_io_in[35]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input31_A (.DIODE(digital_io_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input32_A (.DIODE(digital_io_in[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input33_A (.DIODE(digital_io_in[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input34_A (.DIODE(digital_io_in[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input35_A (.DIODE(digital_io_in[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input36_A (.DIODE(digital_io_in[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input37_A (.DIODE(digital_io_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input38_A (.DIODE(digital_io_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input39_A (.DIODE(e_reset_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input3_A (.DIODE(digital_io_in[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input40_A (.DIODE(i2cm_clk_o));
 sky130_fd_sc_hd__diode_2 ANTENNA_input41_A (.DIODE(i2cm_clk_oen));
 sky130_fd_sc_hd__diode_2 ANTENNA_input42_A (.DIODE(i2cm_data_o));
 sky130_fd_sc_hd__diode_2 ANTENNA_input43_A (.DIODE(i2cm_data_oen));
 sky130_fd_sc_hd__diode_2 ANTENNA_input44_A (.DIODE(i2cm_intr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input45_A (.DIODE(int_pll_clock));
 sky130_fd_sc_hd__diode_2 ANTENNA_input46_A (.DIODE(ir_intr));
 sky130_fd_sc_hd__diode_2 ANTENNA_input47_A (.DIODE(ir_tx));
 sky130_fd_sc_hd__diode_2 ANTENNA_input48_A (.DIODE(p_reset_n));
 sky130_fd_sc_hd__diode_2 ANTENNA_input49_A (.DIODE(reg_addr[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input4_A (.DIODE(digital_io_in[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input50_A (.DIODE(reg_addr[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input51_A (.DIODE(reg_addr[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input52_A (.DIODE(reg_addr[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input53_A (.DIODE(reg_addr[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input54_A (.DIODE(reg_addr[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input55_A (.DIODE(reg_addr[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input56_A (.DIODE(reg_addr[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input57_A (.DIODE(reg_addr[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input58_A (.DIODE(reg_addr[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input59_A (.DIODE(reg_addr[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input5_A (.DIODE(digital_io_in[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input60_A (.DIODE(reg_be[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input61_A (.DIODE(reg_be[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input62_A (.DIODE(reg_be[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input63_A (.DIODE(reg_be[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input64_A (.DIODE(reg_cs));
 sky130_fd_sc_hd__diode_2 ANTENNA_input65_A (.DIODE(reg_peri_ack));
 sky130_fd_sc_hd__diode_2 ANTENNA_input66_A (.DIODE(reg_peri_rdata[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input67_A (.DIODE(reg_peri_rdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input68_A (.DIODE(reg_peri_rdata[11]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input69_A (.DIODE(reg_peri_rdata[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input6_A (.DIODE(digital_io_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input70_A (.DIODE(reg_peri_rdata[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input71_A (.DIODE(reg_peri_rdata[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input72_A (.DIODE(reg_peri_rdata[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input73_A (.DIODE(reg_peri_rdata[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input74_A (.DIODE(reg_peri_rdata[17]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input75_A (.DIODE(reg_peri_rdata[18]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input76_A (.DIODE(reg_peri_rdata[19]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input77_A (.DIODE(reg_peri_rdata[1]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input78_A (.DIODE(reg_peri_rdata[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input79_A (.DIODE(reg_peri_rdata[21]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input7_A (.DIODE(digital_io_in[13]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input80_A (.DIODE(reg_peri_rdata[22]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input81_A (.DIODE(reg_peri_rdata[23]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input82_A (.DIODE(reg_peri_rdata[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input83_A (.DIODE(reg_peri_rdata[25]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input84_A (.DIODE(reg_peri_rdata[26]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input85_A (.DIODE(reg_peri_rdata[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input86_A (.DIODE(reg_peri_rdata[28]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input87_A (.DIODE(reg_peri_rdata[29]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input88_A (.DIODE(reg_peri_rdata[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input89_A (.DIODE(reg_peri_rdata[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input8_A (.DIODE(digital_io_in[14]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input90_A (.DIODE(reg_peri_rdata[31]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input91_A (.DIODE(reg_peri_rdata[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input92_A (.DIODE(reg_peri_rdata[4]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input93_A (.DIODE(reg_peri_rdata[5]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input94_A (.DIODE(reg_peri_rdata[6]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input95_A (.DIODE(reg_peri_rdata[7]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input96_A (.DIODE(reg_peri_rdata[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input97_A (.DIODE(reg_peri_rdata[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input98_A (.DIODE(reg_wdata[0]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input99_A (.DIODE(reg_wdata[10]));
 sky130_fd_sc_hd__diode_2 ANTENNA_input9_A (.DIODE(digital_io_in[15]));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1313_A (.DIODE(net1314));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1322_A (.DIODE(net1321));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1431_A (.DIODE(net1432));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1548_A (.DIODE(net1547));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1558_A (.DIODE(net1557));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length1570_A (.DIODE(net1569));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length5_A (.DIODE(clknet_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_max_length721_A (.DIODE(net720));
 sky130_fd_sc_hd__diode_2 ANTENNA_output199_A (.DIODE(net199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output200_A (.DIODE(net200));
 sky130_fd_sc_hd__diode_2 ANTENNA_output201_A (.DIODE(net201));
 sky130_fd_sc_hd__diode_2 ANTENNA_output202_A (.DIODE(net202));
 sky130_fd_sc_hd__diode_2 ANTENNA_output203_A (.DIODE(net203));
 sky130_fd_sc_hd__diode_2 ANTENNA_output204_A (.DIODE(net204));
 sky130_fd_sc_hd__diode_2 ANTENNA_output205_A (.DIODE(net205));
 sky130_fd_sc_hd__diode_2 ANTENNA_output206_A (.DIODE(net206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output207_A (.DIODE(net207));
 sky130_fd_sc_hd__diode_2 ANTENNA_output208_A (.DIODE(net208));
 sky130_fd_sc_hd__diode_2 ANTENNA_output209_A (.DIODE(net209));
 sky130_fd_sc_hd__diode_2 ANTENNA_output210_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_output211_A (.DIODE(net211));
 sky130_fd_sc_hd__diode_2 ANTENNA_output212_A (.DIODE(net212));
 sky130_fd_sc_hd__diode_2 ANTENNA_output213_A (.DIODE(net213));
 sky130_fd_sc_hd__diode_2 ANTENNA_output214_A (.DIODE(net214));
 sky130_fd_sc_hd__diode_2 ANTENNA_output215_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_output216_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_output217_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_output218_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_output219_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_output220_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_output221_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_output222_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_output223_A (.DIODE(net223));
 sky130_fd_sc_hd__diode_2 ANTENNA_output224_A (.DIODE(net224));
 sky130_fd_sc_hd__diode_2 ANTENNA_output225_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_output226_A (.DIODE(net1108));
 sky130_fd_sc_hd__diode_2 ANTENNA_output227_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_output228_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_output229_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_output230_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_output231_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_output253_A (.DIODE(net253));
 sky130_fd_sc_hd__diode_2 ANTENNA_output254_A (.DIODE(net254));
 sky130_fd_sc_hd__diode_2 ANTENNA_output255_A (.DIODE(net255));
 sky130_fd_sc_hd__diode_2 ANTENNA_output256_A (.DIODE(net256));
 sky130_fd_sc_hd__diode_2 ANTENNA_output257_A (.DIODE(net257));
 sky130_fd_sc_hd__diode_2 ANTENNA_output258_A (.DIODE(net258));
 sky130_fd_sc_hd__diode_2 ANTENNA_output259_A (.DIODE(net581));
 sky130_fd_sc_hd__diode_2 ANTENNA_output260_A (.DIODE(net582));
 sky130_fd_sc_hd__diode_2 ANTENNA_output261_A (.DIODE(net536));
 sky130_fd_sc_hd__diode_2 ANTENNA_output262_A (.DIODE(net537));
 sky130_fd_sc_hd__diode_2 ANTENNA_output263_A (.DIODE(net538));
 sky130_fd_sc_hd__diode_2 ANTENNA_output264_A (.DIODE(net264));
 sky130_fd_sc_hd__diode_2 ANTENNA_output265_A (.DIODE(net583));
 sky130_fd_sc_hd__diode_2 ANTENNA_output266_A (.DIODE(net602));
 sky130_fd_sc_hd__diode_2 ANTENNA_output267_A (.DIODE(net267));
 sky130_fd_sc_hd__diode_2 ANTENNA_output268_A (.DIODE(net268));
 sky130_fd_sc_hd__diode_2 ANTENNA_output269_A (.DIODE(net269));
 sky130_fd_sc_hd__diode_2 ANTENNA_output270_A (.DIODE(net270));
 sky130_fd_sc_hd__diode_2 ANTENNA_output271_A (.DIODE(net271));
 sky130_fd_sc_hd__diode_2 ANTENNA_output272_A (.DIODE(net272));
 sky130_fd_sc_hd__diode_2 ANTENNA_output275_A (.DIODE(net275));
 sky130_fd_sc_hd__diode_2 ANTENNA_output284_A (.DIODE(net284));
 sky130_fd_sc_hd__diode_2 ANTENNA_output285_A (.DIODE(net285));
 sky130_fd_sc_hd__diode_2 ANTENNA_output286_A (.DIODE(net286));
 sky130_fd_sc_hd__diode_2 ANTENNA_output287_A (.DIODE(net287));
 sky130_fd_sc_hd__diode_2 ANTENNA_output288_A (.DIODE(net288));
 sky130_fd_sc_hd__diode_2 ANTENNA_output289_A (.DIODE(net289));
 sky130_fd_sc_hd__diode_2 ANTENNA_output290_A (.DIODE(net290));
 sky130_fd_sc_hd__diode_2 ANTENNA_output291_A (.DIODE(net291));
 sky130_fd_sc_hd__diode_2 ANTENNA_output292_A (.DIODE(net292));
 sky130_fd_sc_hd__diode_2 ANTENNA_output293_A (.DIODE(net293));
 sky130_fd_sc_hd__diode_2 ANTENNA_output294_A (.DIODE(net294));
 sky130_fd_sc_hd__diode_2 ANTENNA_output295_A (.DIODE(net295));
 sky130_fd_sc_hd__diode_2 ANTENNA_output296_A (.DIODE(net529));
 sky130_fd_sc_hd__diode_2 ANTENNA_output297_A (.DIODE(net297));
 sky130_fd_sc_hd__diode_2 ANTENNA_output298_A (.DIODE(net565));
 sky130_fd_sc_hd__diode_2 ANTENNA_output299_A (.DIODE(net530));
 sky130_fd_sc_hd__diode_2 ANTENNA_output300_A (.DIODE(net531));
 sky130_fd_sc_hd__diode_2 ANTENNA_output301_A (.DIODE(net527));
 sky130_fd_sc_hd__diode_2 ANTENNA_output302_A (.DIODE(net302));
 sky130_fd_sc_hd__diode_2 ANTENNA_output303_A (.DIODE(net532));
 sky130_fd_sc_hd__diode_2 ANTENNA_output304_A (.DIODE(net566));
 sky130_fd_sc_hd__diode_2 ANTENNA_output305_A (.DIODE(net305));
 sky130_fd_sc_hd__diode_2 ANTENNA_output306_A (.DIODE(net306));
 sky130_fd_sc_hd__diode_2 ANTENNA_output307_A (.DIODE(net307));
 sky130_fd_sc_hd__diode_2 ANTENNA_output308_A (.DIODE(net308));
 sky130_fd_sc_hd__diode_2 ANTENNA_output309_A (.DIODE(net309));
 sky130_fd_sc_hd__diode_2 ANTENNA_output310_A (.DIODE(net310));
 sky130_fd_sc_hd__diode_2 ANTENNA_output311_A (.DIODE(net1199));
 sky130_fd_sc_hd__diode_2 ANTENNA_output312_A (.DIODE(net1197));
 sky130_fd_sc_hd__diode_2 ANTENNA_output313_A (.DIODE(net313));
 sky130_fd_sc_hd__diode_2 ANTENNA_output314_A (.DIODE(net1195));
 sky130_fd_sc_hd__diode_2 ANTENNA_output315_A (.DIODE(net1193));
 sky130_fd_sc_hd__diode_2 ANTENNA_output316_A (.DIODE(net1191));
 sky130_fd_sc_hd__diode_2 ANTENNA_output317_A (.DIODE(net1189));
 sky130_fd_sc_hd__diode_2 ANTENNA_output318_A (.DIODE(net1187));
 sky130_fd_sc_hd__diode_2 ANTENNA_output319_A (.DIODE(net1185));
 sky130_fd_sc_hd__diode_2 ANTENNA_output320_A (.DIODE(net1183));
 sky130_fd_sc_hd__diode_2 ANTENNA_output321_A (.DIODE(net321));
 sky130_fd_sc_hd__diode_2 ANTENNA_output322_A (.DIODE(net322));
 sky130_fd_sc_hd__diode_2 ANTENNA_output323_A (.DIODE(net323));
 sky130_fd_sc_hd__diode_2 ANTENNA_output324_A (.DIODE(net324));
 sky130_fd_sc_hd__diode_2 ANTENNA_output325_A (.DIODE(net325));
 sky130_fd_sc_hd__diode_2 ANTENNA_output326_A (.DIODE(net528));
 sky130_fd_sc_hd__diode_2 ANTENNA_output327_A (.DIODE(net327));
 sky130_fd_sc_hd__diode_2 ANTENNA_output328_A (.DIODE(net328));
 sky130_fd_sc_hd__diode_2 ANTENNA_output329_A (.DIODE(net329));
 sky130_fd_sc_hd__diode_2 ANTENNA_output330_A (.DIODE(net330));
 sky130_fd_sc_hd__diode_2 ANTENNA_output333_A (.DIODE(net333));
 sky130_fd_sc_hd__diode_2 ANTENNA_output334_A (.DIODE(net334));
 sky130_fd_sc_hd__diode_2 ANTENNA_output335_A (.DIODE(net335));
 sky130_fd_sc_hd__diode_2 ANTENNA_output337_A (.DIODE(net337));
 sky130_fd_sc_hd__diode_2 ANTENNA_output338_A (.DIODE(net338));
 sky130_fd_sc_hd__diode_2 ANTENNA_output339_A (.DIODE(net339));
 sky130_fd_sc_hd__diode_2 ANTENNA_output340_A (.DIODE(net340));
 sky130_fd_sc_hd__diode_2 ANTENNA_output341_A (.DIODE(net341));
 sky130_fd_sc_hd__diode_2 ANTENNA_output342_A (.DIODE(net342));
 sky130_fd_sc_hd__diode_2 ANTENNA_output343_A (.DIODE(net343));
 sky130_fd_sc_hd__diode_2 ANTENNA_output344_A (.DIODE(net344));
 sky130_fd_sc_hd__diode_2 ANTENNA_output345_A (.DIODE(net345));
 sky130_fd_sc_hd__diode_2 ANTENNA_output346_A (.DIODE(net346));
 sky130_fd_sc_hd__diode_2 ANTENNA_output347_A (.DIODE(net347));
 sky130_fd_sc_hd__diode_2 ANTENNA_output348_A (.DIODE(net348));
 sky130_fd_sc_hd__diode_2 ANTENNA_output355_A (.DIODE(net355));
 sky130_fd_sc_hd__diode_2 ANTENNA_output358_A (.DIODE(net358));
 sky130_fd_sc_hd__diode_2 ANTENNA_output359_A (.DIODE(net359));
 sky130_fd_sc_hd__diode_2 ANTENNA_output360_A (.DIODE(net360));
 sky130_fd_sc_hd__diode_2 ANTENNA_output361_A (.DIODE(net361));
 sky130_fd_sc_hd__diode_2 ANTENNA_output362_A (.DIODE(net362));
 sky130_fd_sc_hd__diode_2 ANTENNA_output363_A (.DIODE(net363));
 sky130_fd_sc_hd__diode_2 ANTENNA_output364_A (.DIODE(net364));
 sky130_fd_sc_hd__diode_2 ANTENNA_output365_A (.DIODE(net1206));
 sky130_fd_sc_hd__diode_2 ANTENNA_output366_A (.DIODE(net533));
 sky130_fd_sc_hd__diode_2 ANTENNA_output368_A (.DIODE(net1703));
 sky130_fd_sc_hd__diode_2 ANTENNA_output369_A (.DIODE(net369));
 sky130_fd_sc_hd__diode_2 ANTENNA_output371_A (.DIODE(net371));
 sky130_fd_sc_hd__diode_2 ANTENNA_output373_A (.DIODE(net373));
 sky130_fd_sc_hd__diode_2 ANTENNA_output374_A (.DIODE(net374));
 sky130_fd_sc_hd__diode_2 ANTENNA_output375_A (.DIODE(net375));
 sky130_fd_sc_hd__diode_2 ANTENNA_output376_A (.DIODE(net376));
 sky130_fd_sc_hd__diode_2 ANTENNA_output418_A (.DIODE(net1745));
 sky130_fd_sc_hd__diode_2 ANTENNA_output419_A (.DIODE(net1763));
 sky130_fd_sc_hd__diode_2 ANTENNA_output420_A (.DIODE(net1724));
 sky130_fd_sc_hd__diode_2 ANTENNA_output421_A (.DIODE(net1718));
 sky130_fd_sc_hd__diode_2 ANTENNA_output428_A (.DIODE(net1796));
 sky130_fd_sc_hd__diode_2 ANTENNA_output430_A (.DIODE(net1812));
 sky130_fd_sc_hd__diode_2 ANTENNA_output431_A (.DIODE(net1805));
 sky130_fd_sc_hd__diode_2 ANTENNA_output432_A (.DIODE(net1786));
 sky130_fd_sc_hd__diode_2 ANTENNA_output433_A (.DIODE(net1802));
 sky130_fd_sc_hd__diode_2 ANTENNA_output435_A (.DIODE(net1782));
 sky130_fd_sc_hd__diode_2 ANTENNA_output436_A (.DIODE(net1799));
 sky130_fd_sc_hd__diode_2 ANTENNA_output437_A (.DIODE(net1809));
 sky130_fd_sc_hd__diode_2 ANTENNA_output438_A (.DIODE(net1792));
 sky130_fd_sc_hd__diode_2 ANTENNA_output440_A (.DIODE(net1748));
 sky130_fd_sc_hd__diode_2 ANTENNA_output441_A (.DIODE(net1774));
 sky130_fd_sc_hd__diode_2 ANTENNA_output442_A (.DIODE(net1766));
 sky130_fd_sc_hd__diode_2 ANTENNA_output443_A (.DIODE(net1751));
 sky130_fd_sc_hd__diode_2 ANTENNA_output444_A (.DIODE(net1754));
 sky130_fd_sc_hd__diode_2 ANTENNA_output445_A (.DIODE(net1757));
 sky130_fd_sc_hd__diode_2 ANTENNA_output447_A (.DIODE(net1733));
 sky130_fd_sc_hd__diode_2 ANTENNA_output449_A (.DIODE(net1760));
 sky130_fd_sc_hd__diode_2 ANTENNA_output450_A (.DIODE(net450));
 sky130_fd_sc_hd__diode_2 ANTENNA_output451_A (.DIODE(net451));
 sky130_fd_sc_hd__diode_2 ANTENNA_output452_A (.DIODE(net452));
 sky130_fd_sc_hd__diode_2 ANTENNA_output453_A (.DIODE(net453));
 sky130_fd_sc_hd__diode_2 ANTENNA_output454_A (.DIODE(net1697));
 sky130_fd_sc_hd__diode_2 ANTENNA_output457_A (.DIODE(net457));
 sky130_fd_sc_hd__diode_2 ANTENNA_output459_A (.DIODE(net459));
 sky130_fd_sc_hd__diode_2 ANTENNA_output460_A (.DIODE(net460));
 sky130_fd_sc_hd__diode_2 ANTENNA_output463_A (.DIODE(net463));
 sky130_fd_sc_hd__diode_2 ANTENNA_output465_A (.DIODE(net465));
 sky130_fd_sc_hd__diode_2 ANTENNA_output466_A (.DIODE(net466));
 sky130_fd_sc_hd__diode_2 ANTENNA_output467_A (.DIODE(net467));
 sky130_fd_sc_hd__diode_2 ANTENNA_output468_A (.DIODE(net468));
 sky130_fd_sc_hd__diode_2 ANTENNA_output469_A (.DIODE(net469));
 sky130_fd_sc_hd__diode_2 ANTENNA_output470_A (.DIODE(net470));
 sky130_fd_sc_hd__diode_2 ANTENNA_output471_A (.DIODE(net471));
 sky130_fd_sc_hd__diode_2 ANTENNA_output472_A (.DIODE(net472));
 sky130_fd_sc_hd__diode_2 ANTENNA_output473_A (.DIODE(net473));
 sky130_fd_sc_hd__diode_2 ANTENNA_output474_A (.DIODE(net474));
 sky130_fd_sc_hd__diode_2 ANTENNA_output475_A (.DIODE(net475));
 sky130_fd_sc_hd__diode_2 ANTENNA_output476_A (.DIODE(net476));
 sky130_fd_sc_hd__diode_2 ANTENNA_output477_A (.DIODE(net477));
 sky130_fd_sc_hd__diode_2 ANTENNA_output478_A (.DIODE(net478));
 sky130_fd_sc_hd__diode_2 ANTENNA_output479_A (.DIODE(net479));
 sky130_fd_sc_hd__diode_2 ANTENNA_output480_A (.DIODE(net480));
 sky130_fd_sc_hd__diode_2 ANTENNA_output481_A (.DIODE(net481));
 sky130_fd_sc_hd__diode_2 ANTENNA_output482_A (.DIODE(net482));
 sky130_fd_sc_hd__diode_2 ANTENNA_output484_A (.DIODE(net484));
 sky130_fd_sc_hd__diode_2 ANTENNA_output485_A (.DIODE(net485));
 sky130_fd_sc_hd__diode_2 ANTENNA_output486_A (.DIODE(net486));
 sky130_fd_sc_hd__diode_2 ANTENNA_output487_A (.DIODE(net487));
 sky130_fd_sc_hd__diode_2 ANTENNA_output488_A (.DIODE(net488));
 sky130_fd_sc_hd__diode_2 ANTENNA_output489_A (.DIODE(net489));
 sky130_fd_sc_hd__diode_2 ANTENNA_output490_A (.DIODE(net490));
 sky130_fd_sc_hd__diode_2 ANTENNA_output491_A (.DIODE(net491));
 sky130_fd_sc_hd__diode_2 ANTENNA_output492_A (.DIODE(net492));
 sky130_fd_sc_hd__diode_2 ANTENNA_output493_A (.DIODE(net493));
 sky130_fd_sc_hd__diode_2 ANTENNA_output494_A (.DIODE(net494));
 sky130_fd_sc_hd__diode_2 ANTENNA_output495_A (.DIODE(net495));
 sky130_fd_sc_hd__diode_2 ANTENNA_output496_A (.DIODE(net496));
 sky130_fd_sc_hd__diode_2 ANTENNA_output502_A (.DIODE(net502));
 sky130_fd_sc_hd__diode_2 ANTENNA_output505_A (.DIODE(net601));
 sky130_fd_sc_hd__diode_2 ANTENNA_output506_A (.DIODE(net506));
 sky130_fd_sc_hd__diode_2 ANTENNA_output509_A (.DIODE(net509));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_cpu0_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[8] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_cpu1_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[9] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_cpu2_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[10] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_cpu3_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[11] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_cpu_intf_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[0] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_i2cm_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[4] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_sspim_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[2] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_uart0_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[3] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_uart1_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[6] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_buf_usb_rst.u_buf_A  (.DIODE(\u_glbl_reg.cfg_rst_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_clkbuf_dbg_ref.u_buf_A  (.DIODE(net1693));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_rtc_clk_sel.genblk1.u_mux_S  (.DIODE(\u_glbl_reg.cfg_rtc_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_glbl_reg.u_usb_clk_sel.genblk1.u_mux_S  (.DIODE(\u_glbl_reg.cfg_usb_clk_ctrl[5] ));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_00.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_01.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_02.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_03.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_04.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_05.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_06.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_07.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_10.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_11.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_12.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_13.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_20.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_21.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[2]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_skew_pinmux.u_mux_level_30.genblk1.u_mux_S  (.DIODE(cfg_cska_pinmux[3]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1043_A (.DIODE(net1042));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1093_A (.DIODE(net222));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1094_A (.DIODE(net221));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1095_A (.DIODE(net220));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1096_A (.DIODE(net219));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1097_A (.DIODE(net218));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1098_A (.DIODE(net217));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1099_A (.DIODE(net210));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1100_A (.DIODE(net225));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1101_A (.DIODE(net231));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1102_A (.DIODE(net230));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1103_A (.DIODE(net229));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1104_A (.DIODE(net228));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1105_A (.DIODE(net227));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1106_A (.DIODE(net216));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1107_A (.DIODE(net215));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1108_A (.DIODE(net226));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1183_A (.DIODE(net1184));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1184_A (.DIODE(net320));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1185_A (.DIODE(net1186));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1186_A (.DIODE(net319));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1187_A (.DIODE(net1188));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1188_A (.DIODE(net318));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1189_A (.DIODE(net1190));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1190_A (.DIODE(net317));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1191_A (.DIODE(net1192));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1192_A (.DIODE(net316));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1193_A (.DIODE(net1194));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1194_A (.DIODE(net315));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1195_A (.DIODE(net1196));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1196_A (.DIODE(net314));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1197_A (.DIODE(net1198));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1198_A (.DIODE(net312));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1199_A (.DIODE(net1200));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1200_A (.DIODE(net311));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1206_A (.DIODE(net365));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1285_A (.DIODE(net1284));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1304_A (.DIODE(net9));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1305_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1306_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1315_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1318_A (.DIODE(net1317));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1386_A (.DIODE(net1385));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1389_A (.DIODE(net1390));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1391_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1393_A (.DIODE(net1394));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1394_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1395_A (.DIODE(net1396));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1396_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1400_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1401_A (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1403_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1404_A (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1406_A (.DIODE(net1407));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1407_A (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1408_A (.DIODE(net1409));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1409_A (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1410_A (.DIODE(net1411));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1411_A (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1412_A (.DIODE(net1413));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1413_A (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1414_A (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1415_A (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1416_A (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1417_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1439_A (.DIODE(net1438));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1455_A (.DIODE(net1454));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1480_A (.DIODE(net1479));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1487_A (.DIODE(net1486));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1495_A (.DIODE(net1494));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1497_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1511_A (.DIODE(net1510));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1518_A (.DIODE(net1517));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1525_A (.DIODE(net1524));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1532_A (.DIODE(net1533));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1540_A (.DIODE(net1539));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1571_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1578_A (.DIODE(net1577));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1588_A (.DIODE(net1587));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1593_A (.DIODE(net1592));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1594_A (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1596_A (.DIODE(net1595));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1605_A (.DIODE(net1604));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1627_A (.DIODE(net1626));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1634_A (.DIODE(net1635));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1642_A (.DIODE(net1641));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1649_A (.DIODE(net1648));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1650_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1652_A (.DIODE(net1651));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1653_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_A (.DIODE(net1694));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire4_A (.DIODE(\u_glbl_reg.dbg_clk_ref ));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire527_A (.DIODE(net301));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire528_A (.DIODE(net326));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire530_A (.DIODE(net299));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire531_A (.DIODE(net300));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire532_A (.DIODE(net303));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire536_A (.DIODE(net261));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire537_A (.DIODE(net262));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire538_A (.DIODE(net263));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire565_A (.DIODE(net298));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire566_A (.DIODE(net304));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire581_A (.DIODE(net259));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire582_A (.DIODE(net260));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire583_A (.DIODE(net265));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire602_A (.DIODE(net266));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire6_A (.DIODE(clknet_0_mclk));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire7_A (.DIODE(net1698));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(net1699));
 sky130_fd_sc_hd__decap_4 FILLER_0_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1029 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1055 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1070 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_560 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_100_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_100_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_100_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_100_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_100_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_100_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_100_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_588 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_666 ();
 sky130_fd_sc_hd__decap_3 FILLER_101_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_712 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_766 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_101_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_101_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_101_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_101_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_101_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_101_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_102_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_102_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_731 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_854 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_102_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_102_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_102_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_102_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_102_992 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_151 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_512 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_103_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_804 ();
 sky130_fd_sc_hd__decap_6 FILLER_103_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_103_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_103_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_103_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_103_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_103_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_1003 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_104_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_270 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_658 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_831 ();
 sky130_fd_sc_hd__decap_8 FILLER_104_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_104_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_104_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_104_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_104_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_104_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_1077 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_26 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_654 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_795 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_801 ();
 sky130_ef_sc_hd__decap_12 FILLER_105_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_105_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_105_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_105_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_105_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_105_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_105_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_106_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1091 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_572 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_106_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_106_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_106_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_106_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_106_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_106_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_1019 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_1089 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_548 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_107_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_828 ();
 sky130_fd_sc_hd__decap_3 FILLER_107_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_107_902 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_107_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_107_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_107_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_107_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1022 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_108_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_571 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_574 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_108_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_108_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_108_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_108_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_108_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_108_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_109_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_256 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_32 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_370 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_109_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_109_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_883 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_109_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_109_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_109_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_109_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_574 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_790 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_800 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_876 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_110_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_794 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_110_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_110_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_110_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_110_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_110_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_110_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1026 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_111_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_111_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_111_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_111_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_111_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_111_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_111_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_1003 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1011 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_112_840 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_112_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_112_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_112_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_112_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_112_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_112_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_862 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_113_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_113_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_113_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_113_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_113_971 ();
 sky130_fd_sc_hd__decap_8 FILLER_113_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1005 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1024 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1064 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_1076 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_218 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_235 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_114_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_616 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_114_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_114_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_114_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_114_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_114_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_114_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1001 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_519 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_578 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_115_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_115_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_115_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_115_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_115_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_115_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_115_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1044 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_116_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_116_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_116_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_116_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_116_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_116_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_116_999 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1018 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_117_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_117_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_117_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_117_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_117_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_117_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_117_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1019 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_1082 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_691 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_900 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_118_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_118_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_118_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_118_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_118_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_118_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_118_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1034 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_1094 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_244 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_580 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_119_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_119_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_119_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_119_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_119_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_119_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_119_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_291 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_668 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_719 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1021 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_1074 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1086 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_454 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_120_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_888 ();
 sky130_ef_sc_hd__decap_12 FILLER_120_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_120_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_120_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_120_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_120_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_120_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1026 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1032 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1042 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_574 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_656 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_121_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_863 ();
 sky130_ef_sc_hd__decap_12 FILLER_121_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_121_887 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_121_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_121_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_121_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_121_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1016 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_180 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_294 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_122_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_122_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_122_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_122_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_122_976 ();
 sky130_fd_sc_hd__decap_3 FILLER_122_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_122_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_123_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_123_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_868 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_123_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_123_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_123_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_123_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_123_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1046 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_1070 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_274 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_124_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_124_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_124_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_124_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_124_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_124_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_124_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_1005 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_125_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_125_837 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_125_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_125_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_125_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_125_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_125_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1014 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_126_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_13 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_835 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_126_948 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_126_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_126_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_126_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_126_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_127_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_144 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_255 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_663 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_127_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_836 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_87 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_127_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_127_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_127_983 ();
 sky130_fd_sc_hd__fill_1 FILLER_127_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_127_998 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1045 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_128_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_128_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_842 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_128_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_128_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_128_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_128_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_128_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1038 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_129_1071 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_129_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_129_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_129_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_129_962 ();
 sky130_fd_sc_hd__decap_8 FILLER_129_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_129_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_598 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_730 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_790 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1014 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1018 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1064 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1073 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_130_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_899 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_130_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_130_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_130_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_130_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_130_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_130_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1006 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1028 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_1035 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1060 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_1072 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_1091 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_13 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_254 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_327 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_782 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_131_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_131_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_131_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_946 ();
 sky130_fd_sc_hd__decap_6 FILLER_131_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_131_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_131_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_131_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_1074 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1082 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_434 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_674 ();
 sky130_fd_sc_hd__decap_6 FILLER_132_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_132_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_837 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_132_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_132_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_132_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_132_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_132_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1029 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1041 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_700 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_816 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_133_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_133_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_920 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_940 ();
 sky130_fd_sc_hd__decap_8 FILLER_133_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_133_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_133_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_133_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_133_992 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_1005 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1032 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_1067 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_776 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_844 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_855 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_134_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_134_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_134_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_134_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_134_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_134_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_134_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1003 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1031 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_258 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_579 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_759 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_864 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_135_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_135_895 ();
 sky130_fd_sc_hd__decap_3 FILLER_135_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_135_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_135_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_135_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_135_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_101 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_282 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_336 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_450 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_136_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_136_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_136_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_136_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_136_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_136_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_136_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1004 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1027 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1033 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1052 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_137_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_137_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_137_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_137_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_137_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_137_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_137_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_1087 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_138_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_138_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_138_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_138_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_138_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_138_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_138_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_364 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_139_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_812 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_139_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_928 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_139_940 ();
 sky130_fd_sc_hd__fill_2 FILLER_139_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_139_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_139_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_139_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_463 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_1097 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_484 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_140_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_140_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_140_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_140_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_140_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_140_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_140_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1087 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_42 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_547 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_141_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_141_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_141_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_141_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_141_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_141_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_141_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_142_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_142_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_142_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_945 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_142_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_142_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_142_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_142_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_1065 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_1088 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_256 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_358 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_378 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_707 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_880 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_884 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_143_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_143_932 ();
 sky130_fd_sc_hd__decap_3 FILLER_143_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_143_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_143_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_143_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_143_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_50 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_144_888 ();
 sky130_fd_sc_hd__fill_1 FILLER_144_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_144_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_144_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_144_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_144_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_144_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_247 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_366 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_145_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_702 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_145_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_145_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_145_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_145_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_145_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_145_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_338 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_578 ();
 sky130_fd_sc_hd__decap_3 FILLER_146_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_146_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_146_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_146_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_146_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_146_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_146_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_666 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_819 ();
 sky130_fd_sc_hd__decap_6 FILLER_147_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_147_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_147_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_917 ();
 sky130_fd_sc_hd__decap_3 FILLER_147_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_147_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_147_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_147_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_228 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_432 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_602 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_148_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_148_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_148_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_148_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_148_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_148_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_148_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_149_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_149_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_882 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_149_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_149_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_149_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_149_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_149_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_227 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_619 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_1073 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_1085 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_562 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_150_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_150_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_150_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_150_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_150_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_150_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_150_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_1077 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_151_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_586 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_833 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_151_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_151_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_151_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_151_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_151_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_151_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_14 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_152_711 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_731 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_152_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_152_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_901 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_152_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_152_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_152_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_152_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_243 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_36 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_430 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_153_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_153_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_153_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_940 ();
 sky130_fd_sc_hd__decap_6 FILLER_153_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_153_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_153_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_153_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_170 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_284 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_842 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_154_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_154_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_154_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_154_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_154_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_154_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_154_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_10 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_198 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_155_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_155_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_155_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_155_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_957 ();
 sky130_fd_sc_hd__decap_3 FILLER_155_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_155_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_155_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_901 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_156_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_156_941 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_156_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_156_978 ();
 sky130_fd_sc_hd__decap_8 FILLER_156_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_156_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_156_992 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_744 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_157_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_157_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_157_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_933 ();
 sky130_fd_sc_hd__fill_1 FILLER_157_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_157_940 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_953 ();
 sky130_fd_sc_hd__decap_3 FILLER_157_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_157_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_665 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_735 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_158_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_158_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_158_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_158_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_158_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_158_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_158_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_159_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_159_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_159_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_159_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_159_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_159_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_159_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_597 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_644 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_845 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_977 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_507 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_8 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_160_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_160_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_920 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_160_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_160_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_160_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_160_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_160_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_161_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_681 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_161_927 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_936 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_161_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_161_963 ();
 sky130_fd_sc_hd__fill_2 FILLER_161_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_161_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_161_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_302 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_344 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_861 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_162_918 ();
 sky130_fd_sc_hd__decap_3 FILLER_162_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_162_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_162_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_162_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_162_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_162_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_163_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_163_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_163_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_163_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_163_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_163_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_163_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_1093 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_213 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_290 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_605 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_164_898 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_164_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_164_931 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_164_957 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_164_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_164_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_164_996 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_165_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_903 ();
 sky130_fd_sc_hd__decap_6 FILLER_165_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_165_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_165_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_165_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_165_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_165_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_166_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_166_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_789 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_166_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_898 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_166_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_166_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_166_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_166_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_1058 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_167_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_167_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_527 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_592 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_703 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_710 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_167_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_167_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_167_963 ();
 sky130_fd_sc_hd__decap_6 FILLER_167_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_167_997 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1034 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1084 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_548 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_168_823 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_168_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_168_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_168_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_168_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_168_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_168_981 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1009 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_1043 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_659 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_808 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_169_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_169_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_169_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_169_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_169_987 ();
 sky130_fd_sc_hd__fill_1 FILLER_169_995 ();
 sky130_fd_sc_hd__decap_4 FILLER_169_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_342 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_376 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_730 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1014 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_1025 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1034 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1043 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1055 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1067 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_1079 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_555 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_572 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_170_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_835 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_170_903 ();
 sky130_fd_sc_hd__decap_3 FILLER_170_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_170_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_170_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_170_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_170_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_407 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_580 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_818 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_171_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_171_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_171_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_171_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_171_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_171_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_171_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_1003 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1015 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1021 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_715 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_172_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_172_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_172_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_172_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_172_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_172_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_172_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_173_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_28 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_429 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_465 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_768 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_173_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_870 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_173_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_173_953 ();
 sky130_fd_sc_hd__decap_8 FILLER_173_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_173_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_173_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_483 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_174_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_174_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_852 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_174_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_174_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_174_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_174_981 ();
 sky130_fd_sc_hd__decap_8 FILLER_174_985 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1015 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_367 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_175_797 ();
 sky130_fd_sc_hd__decap_6 FILLER_175_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_175_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_175_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_175_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_175_986 ();
 sky130_fd_sc_hd__decap_4 FILLER_175_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_804 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_833 ();
 sky130_fd_sc_hd__decap_8 FILLER_176_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_176_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_176_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_176_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_176_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_176_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_176_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_1056 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_371 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_482 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_772 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_816 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_828 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_177_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_177_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_177_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_177_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_177_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_177_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_177_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_1017 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_124 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_750 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_781 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_178_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_178_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_178_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_178_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_178_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_178_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_178_995 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1031 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1039 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_146 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_252 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_179_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_179_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_179_937 ();
 sky130_fd_sc_hd__fill_2 FILLER_179_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_179_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_976 ();
 sky130_fd_sc_hd__decap_4 FILLER_179_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_179_988 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_256 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_368 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_714 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_720 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_865 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_877 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_17_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_1030 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1045 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1057 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_1069 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1081 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_1089 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_491 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_180_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_891 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_180_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_180_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_180_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_180_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_180_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_180_991 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_1017 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_161 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_194 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_267 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_710 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_181_766 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_792 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_824 ();
 sky130_fd_sc_hd__decap_3 FILLER_181_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_181_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_181_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_181_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_181_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_181_996 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1004 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_1012 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1020 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_549 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_182_921 ();
 sky130_fd_sc_hd__decap_6 FILLER_182_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_182_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_182_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_182_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_182_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_182_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_1021 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1046 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_1058 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_31 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_319 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_422 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_812 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_818 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_863 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_870 ();
 sky130_fd_sc_hd__fill_1 FILLER_183_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_886 ();
 sky130_fd_sc_hd__decap_6 FILLER_183_89 ();
 sky130_fd_sc_hd__decap_3 FILLER_183_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_916 ();
 sky130_fd_sc_hd__decap_8 FILLER_183_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_183_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_183_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_183_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_172 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_210 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_435 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_664 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_184_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_921 ();
 sky130_fd_sc_hd__decap_3 FILLER_184_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_184_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_184_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_184_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_184_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_184_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_192 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_426 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_812 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_857 ();
 sky130_fd_sc_hd__decap_8 FILLER_185_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_890 ();
 sky130_fd_sc_hd__decap_3 FILLER_185_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_915 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_185_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_185_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_185_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_185_969 ();
 sky130_fd_sc_hd__fill_2 FILLER_185_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_186_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_148 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_158 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_563 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_186_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_186_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_806 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_186_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_186_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_186_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_186_996 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_1018 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1027 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1039 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1051 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_520 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_542 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_637 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_187_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_814 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_826 ();
 sky130_fd_sc_hd__decap_3 FILLER_187_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_187_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_187_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_187_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_187_975 ();
 sky130_fd_sc_hd__decap_8 FILLER_187_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1013 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_188_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_188_757 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_188_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_188_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_188_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_188_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_188_990 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_1013 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_1020 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_371 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_189_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_189_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_189_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_189_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_189_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_189_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_189_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_571 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_836 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_906 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_101 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1011 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_25 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_190_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_190_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_190_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_190_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_190_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_190_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_190_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1000 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_1023 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1042 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_1054 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1062 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_772 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_191_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_888 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_191_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_915 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_939 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_191_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_191_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_191_975 ();
 sky130_fd_sc_hd__decap_3 FILLER_191_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_191_988 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1004 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_130 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_262 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_283 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_352 ();
 sky130_fd_sc_hd__decap_3 FILLER_192_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_192_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_776 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_192_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_192_976 ();
 sky130_fd_sc_hd__decap_6 FILLER_192_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_192_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_192_992 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1022 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1036 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1048 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_471 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_600 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_606 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_193_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_807 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_872 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_193_906 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_193_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_193_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_193_98 ();
 sky130_fd_sc_hd__decap_3 FILLER_193_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_193_996 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1010 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_14 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_46 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_59 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_843 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_194_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_194_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_194_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_194_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_194_959 ();
 sky130_fd_sc_hd__decap_3 FILLER_194_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_194_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_1002 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_1055 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_420 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_195_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_752 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_195_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_851 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_195_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_195_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_195_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_195_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_195_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_196_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_490 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_594 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_8 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_196_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_196_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_196_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_96 ();
 sky130_fd_sc_hd__decap_4 FILLER_196_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_196_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_196_994 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_1002 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1029 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1041 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_1053 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_176 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_25 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_606 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_197_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_197_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_197_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_197_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_197_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_960 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_966 ();
 sky130_ef_sc_hd__decap_12 FILLER_197_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_197_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_292 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_675 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_684 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_198_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_198_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_198_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_198_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_198_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_981 ();
 sky130_fd_sc_hd__decap_6 FILLER_198_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_198_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_132 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_20 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_199_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_199_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_199_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_199_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_199_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_199_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_199_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_439 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_606 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_804 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1038 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1044 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1050 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1058 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1062 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_18 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_415 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_427 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_54 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_36 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_608 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_786 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_200_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_200_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_200_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_200_944 ();
 sky130_fd_sc_hd__decap_4 FILLER_200_95 ();
 sky130_fd_sc_hd__decap_8 FILLER_200_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_200_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_10 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_22 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_361 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_201_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_201_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_201_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_201_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_201_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_201_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_201_988 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_324 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_450 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_46 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_564 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_632 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_695 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_749 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_829 ();
 sky130_fd_sc_hd__decap_6 FILLER_202_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_202_862 ();
 sky130_fd_sc_hd__decap_3 FILLER_202_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_929 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_202_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_958 ();
 sky130_fd_sc_hd__decap_8 FILLER_202_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_202_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_202_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_500 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_203_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_650 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_203_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_789 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_203_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_203_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_203_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_203_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_203_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_216 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_38 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_439 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_204_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_607 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_636 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_788 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_792 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_204_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_204_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_921 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_204_933 ();
 sky130_fd_sc_hd__decap_8 FILLER_204_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_204_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_204_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_199 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_384 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_488 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_205_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_801 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_205_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_205_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_205_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_205_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_205_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_205_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_168 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_444 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_206_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_50 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_206_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_538 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_790 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_798 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_206_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_206_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_206_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_206_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_206_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_260 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_471 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_514 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_207_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_207_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_207_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_873 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_207_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_207_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_207_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_207_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_115 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_493 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_597 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_682 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_208_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_208_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_208_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_208_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_208_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_208_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_208_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1045 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_120 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_19 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_198 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_232 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_303 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_311 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_209_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_882 ();
 sky130_fd_sc_hd__decap_3 FILLER_209_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_915 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_209_938 ();
 sky130_fd_sc_hd__fill_1 FILLER_209_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_209_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_209_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_968 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_980 ();
 sky130_ef_sc_hd__decap_12 FILLER_209_992 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_654 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_56 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_723 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_762 ();
 sky130_fd_sc_hd__decap_8 FILLER_210_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_795 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_210_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_210_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_210_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_210_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_962 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_210_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_210_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_693 ();
 sky130_fd_sc_hd__decap_3 FILLER_211_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_756 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_814 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_820 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_211_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_211_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_211_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_211_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_211_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_211_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_189 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_212_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_623 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_735 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_212_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_900 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_912 ();
 sky130_fd_sc_hd__decap_8 FILLER_212_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_212_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_212_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_212_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_212_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_270 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_213_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_841 ();
 sky130_fd_sc_hd__decap_3 FILLER_213_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_213_930 ();
 sky130_fd_sc_hd__fill_2 FILLER_213_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_213_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_213_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_213_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1029 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_146 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_38 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_400 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_486 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_214_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_214_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_891 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_214_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_214_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_214_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_214_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_214_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_458 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_464 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_215_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_215_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_215_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_215_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_215_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_215_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_215_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1017 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_36 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_216_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_681 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_216_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_216_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_216_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_957 ();
 sky130_fd_sc_hd__decap_8 FILLER_216_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_216_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_216_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1045 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_191 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_269 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_31 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_404 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_422 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_217_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_217_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_217_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_217_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_217_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_965 ();
 sky130_fd_sc_hd__decap_8 FILLER_217_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_217_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_1085 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_241 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_247 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_427 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_448 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_486 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_578 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_218_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_218_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_667 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_689 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_218_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_875 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_218_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_218_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_218_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_218_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_245 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_523 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_691 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_219_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_825 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_219_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_219_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_219_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_219_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_219_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_219_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_639 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_642 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_749 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_760 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_808 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_853 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_865 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_562 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_674 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_697 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_220_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_728 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_785 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_220_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_220_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_220_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_220_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_220_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_220_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_267 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_376 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_550 ();
 sky130_fd_sc_hd__decap_3 FILLER_221_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_221_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_221_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_876 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_221_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_221_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_221_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_221_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_118 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_734 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_222_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_874 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_222_904 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_222_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_222_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_222_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_222_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_222_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_406 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_456 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_656 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_758 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_839 ();
 sky130_fd_sc_hd__decap_3 FILLER_223_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_223_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_223_921 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_223_934 ();
 sky130_fd_sc_hd__decap_8 FILLER_223_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_223_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_223_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_275 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_388 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_490 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_611 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_224_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_224_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_224_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_224_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_224_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_224_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_224_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_372 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_480 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_600 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_636 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_739 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_225_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_225_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_225_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_225_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_225_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_225_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_225_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_226_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_226_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_840 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_874 ();
 sky130_fd_sc_hd__fill_1 FILLER_226_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_226_964 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_226_970 ();
 sky130_fd_sc_hd__fill_2 FILLER_226_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_226_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_142 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_479 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_801 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_821 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_227_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_859 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_227_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_227_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_227_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_227_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_227_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_227_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_683 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_778 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_799 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_842 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_228_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_228_886 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_228_925 ();
 sky130_fd_sc_hd__fill_2 FILLER_228_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_228_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_228_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_228_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_298 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_418 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_792 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_845 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_229_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_229_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_229_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_911 ();
 sky130_fd_sc_hd__decap_8 FILLER_229_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_229_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_229_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_229_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_216 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_331 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_878 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_229 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_230_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_828 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_834 ();
 sky130_fd_sc_hd__decap_6 FILLER_230_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_230_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_230_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_939 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_230_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_230_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_230_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_127 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_216 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_420 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_540 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_231_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_766 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_815 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_819 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_231_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_231_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_231_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_231_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_231_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_231_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_204 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_212 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_402 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_609 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_654 ();
 sky130_fd_sc_hd__decap_3 FILLER_232_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_685 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_774 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_787 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_832 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_885 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_232_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_232_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_232_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_232_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_232_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_232_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1033 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_288 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_350 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_233_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_708 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_714 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_863 ();
 sky130_fd_sc_hd__decap_8 FILLER_233_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_233_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_233_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_233_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_233_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_233_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_512 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_555 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_234_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_234_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_873 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_234_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_234_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_234_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_234_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_234_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_427 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_235_696 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_716 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_235_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_867 ();
 sky130_fd_sc_hd__fill_1 FILLER_235_871 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_235_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_235_919 ();
 sky130_fd_sc_hd__fill_2 FILLER_235_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_235_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_243 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_707 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_236_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_823 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_860 ();
 sky130_fd_sc_hd__decap_3 FILLER_236_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_910 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_236_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_236_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_236_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_236_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_236_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_1057 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_182 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_268 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_476 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_783 ();
 sky130_fd_sc_hd__decap_6 FILLER_237_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_793 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_818 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_853 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_237_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_911 ();
 sky130_fd_sc_hd__decap_3 FILLER_237_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_237_932 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_938 ();
 sky130_fd_sc_hd__fill_2 FILLER_237_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_977 ();
 sky130_fd_sc_hd__decap_8 FILLER_237_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_237_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_584 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_74 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_788 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_238_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_238_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_238_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_238_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_238_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_238_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_238_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_140 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_315 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_440 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_488 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_239_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_758 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_239_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_239_808 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_847 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_239_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_239_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_239_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_239_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_198 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_583 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_595 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_722 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_742 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_23_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_917 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_236 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_507 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_240_843 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_881 ();
 sky130_fd_sc_hd__decap_6 FILLER_240_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_905 ();
 sky130_fd_sc_hd__decap_8 FILLER_240_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_240_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_240_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_240_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_240_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_1089 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_426 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_241_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_241_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_241_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_241_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_241_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_241_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_241_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_406 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_242_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_846 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_242_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_242_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_887 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_242_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_242_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_242_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_242_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_412 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_462 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_243_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_243_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_854 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_884 ();
 sky130_fd_sc_hd__decap_8 FILLER_243_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_243_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_243_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_243_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_243_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_544 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_720 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_740 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_858 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_244_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_244_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_914 ();
 sky130_fd_sc_hd__decap_3 FILLER_244_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_244_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_244_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_244_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_244_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_290 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_494 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_510 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_781 ();
 sky130_fd_sc_hd__decap_8 FILLER_245_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_793 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_798 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_245_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_245_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_245_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_245_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_245_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_245_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_575 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_59 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_634 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_767 ();
 sky130_fd_sc_hd__decap_3 FILLER_246_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_784 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_840 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_880 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_246_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_246_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_246_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_246_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_246_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_246_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_359 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_485 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_573 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_745 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_798 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_247_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_247_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_902 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_247_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_247_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_247_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_247_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_247_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_117 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_369 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_405 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_696 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_248_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_248_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_248_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_907 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_248_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_248_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_248_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_248_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_308 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_404 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_518 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_688 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_715 ();
 sky130_fd_sc_hd__decap_3 FILLER_249_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_780 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_807 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_249_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_249_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_249_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_249_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_249_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_249_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_269 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_58 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_734 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_851 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_898 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_23 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_443 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_603 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_619 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_250_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_731 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_250_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_802 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_250_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_250_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_250_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_250_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_250_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_218 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_255 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_476 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_482 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_67 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_251_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_251_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_850 ();
 sky130_fd_sc_hd__decap_8 FILLER_251_860 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_878 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_251_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_251_926 ();
 sky130_fd_sc_hd__fill_2 FILLER_251_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_251_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_151 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_243 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_392 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_510 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_571 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_674 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_736 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_783 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_824 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_830 ();
 sky130_fd_sc_hd__decap_3 FILLER_252_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_252_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_252_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_252_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_252_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_252_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_252_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_144 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_478 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_491 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_253_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_597 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_253_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_803 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_253_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_253_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_253_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_253_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_253_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_496 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_508 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_679 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_827 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_846 ();
 sky130_fd_sc_hd__decap_3 FILLER_254_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_254_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_878 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_254_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_254_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_254_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_254_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_254_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_472 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_689 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_706 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_795 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_255_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_255_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_846 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_255_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_255_945 ();
 sky130_fd_sc_hd__decap_8 FILLER_255_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_255_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_255_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_151 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_256_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_708 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_722 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_836 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_857 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_256_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_256_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_256_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_256_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_256_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_256_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_257_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_549 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_257_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_257_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_257_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_257_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_257_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_257_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1005 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_1085 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_272 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_455 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_551 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_668 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_672 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_735 ();
 sky130_fd_sc_hd__decap_3 FILLER_258_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_781 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_787 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_796 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_877 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_258_910 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_258_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_258_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_258_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_962 ();
 sky130_fd_sc_hd__decap_6 FILLER_258_974 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_258_993 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_160 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_238 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_329 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_411 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_700 ();
 sky130_fd_sc_hd__decap_3 FILLER_259_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_862 ();
 sky130_fd_sc_hd__decap_8 FILLER_259_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_259_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_259_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_259_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_259_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_958 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_970 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_982 ();
 sky130_ef_sc_hd__decap_12 FILLER_259_994 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_43 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_594 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_607 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_755 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_882 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_121 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_163 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_260_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_430 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_260_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_260_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_873 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_885 ();
 sky130_fd_sc_hd__decap_8 FILLER_260_908 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_260_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_956 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_260_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_260_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_372 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_403 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_609 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_850 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_261_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_872 ();
 sky130_fd_sc_hd__decap_8 FILLER_261_881 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_889 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_261_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_261_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_261_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_261_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_261_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_412 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_547 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_262_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_818 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_831 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_849 ();
 sky130_fd_sc_hd__decap_6 FILLER_262_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_852 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_905 ();
 sky130_fd_sc_hd__fill_1 FILLER_262_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_262_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_262_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_262_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_262_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_368 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_408 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_480 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_567 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_759 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_826 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_263_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_847 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_86 ();
 sky130_fd_sc_hd__decap_3 FILLER_263_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_880 ();
 sky130_fd_sc_hd__decap_6 FILLER_263_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_263_895 ();
 sky130_fd_sc_hd__decap_8 FILLER_263_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_263_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_263_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_126 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_154 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_676 ();
 sky130_fd_sc_hd__decap_6 FILLER_264_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_727 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_786 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_792 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_264_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_264_824 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_891 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_264_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_264_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_264_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_264_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_399 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_442 ();
 sky130_fd_sc_hd__decap_3 FILLER_265_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_591 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_630 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_758 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_265_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_265_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_870 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_909 ();
 sky130_fd_sc_hd__decap_6 FILLER_265_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_265_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_265_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_265_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_340 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_772 ();
 sky130_fd_sc_hd__decap_8 FILLER_266_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_788 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_266_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_840 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_876 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_900 ();
 sky130_fd_sc_hd__fill_2 FILLER_266_922 ();
 sky130_fd_sc_hd__decap_3 FILLER_266_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_933 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_952 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_964 ();
 sky130_fd_sc_hd__decap_6 FILLER_266_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_266_976 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_266_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_262 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_316 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_328 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_454 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_535 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_598 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_639 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_267_789 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_824 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_267_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_267_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_267_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_267_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_267_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_267_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_192 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_441 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_751 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_268_876 ();
 sky130_fd_sc_hd__decap_6 FILLER_268_884 ();
 sky130_fd_sc_hd__fill_1 FILLER_268_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_268_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_909 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_917 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_268_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_268_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_268_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_269_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_269_669 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_804 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_832 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_269_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_269_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_916 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_269_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_269_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_269_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_260 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_340 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_360 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_370 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_712 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_883 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1017 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_122 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_175 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_270_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_623 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_270_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_854 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_270_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_270_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_270_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_270_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_270_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_348 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_271_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_768 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_807 ();
 sky130_fd_sc_hd__decap_3 FILLER_271_815 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_870 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_904 ();
 sky130_fd_sc_hd__decap_6 FILLER_271_913 ();
 sky130_fd_sc_hd__decap_8 FILLER_271_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_271_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_271_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_271_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_179 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_339 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_466 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_624 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_744 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_77 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_784 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_830 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_849 ();
 sky130_fd_sc_hd__decap_3 FILLER_272_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_272_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_272_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_910 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_272_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_272_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_936 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_948 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_960 ();
 sky130_fd_sc_hd__decap_8 FILLER_272_972 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_272_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_202 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_600 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_826 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_273_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_861 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_873 ();
 sky130_fd_sc_hd__decap_8 FILLER_273_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_273_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_273_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_273_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_905 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_273_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_273_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_1085 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_13 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_315 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_353 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_512 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_681 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_717 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_274_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_806 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_274_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_274_893 ();
 sky130_fd_sc_hd__decap_3 FILLER_274_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_274_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_274_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_274_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_11 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_352 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_479 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_635 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_733 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_275_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_275_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_275_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_845 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_275_860 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_275_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_275_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_275_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_735 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_276_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_276_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_848 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_890 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_276_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_276_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_276_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_276_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_276_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_17 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_300 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_319 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_375 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_550 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_727 ();
 sky130_fd_sc_hd__decap_3 FILLER_277_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_796 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_808 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_277_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_877 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_277_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_277_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_277_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_277_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_277_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_34 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_418 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_444 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_560 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_572 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_278_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_719 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_732 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_796 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_278_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_278_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_278_915 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_278_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_278_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_278_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_16 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_355 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_367 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_715 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_279_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_279_775 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_808 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_279_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_279_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_279_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_913 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_279_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_279_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_38 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_603 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_780 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_893 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_926 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_68 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_280_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_776 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_800 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_280_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_867 ();
 sky130_fd_sc_hd__decap_3 FILLER_280_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_280_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_280_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_280_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_280_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_816 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_822 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_281_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_281_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_858 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_281_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_281_937 ();
 sky130_fd_sc_hd__decap_8 FILLER_281_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_281_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_281_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_214 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_339 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_409 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_523 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_600 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_734 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_282_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_824 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_859 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_282_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_282_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_282_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_282_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_282_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_282_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_22 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_312 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_325 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_511 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_628 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_640 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_646 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_283_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_283_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_283_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_927 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_283_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_283_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_283_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_969 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_283_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1005 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_14 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_474 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_643 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_284_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_284_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_284_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_284_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_957 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_284_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_284_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_284_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_1101 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_418 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_285_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_637 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_687 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_775 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_827 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_830 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_838 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_880 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_285_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_285_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_285_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_285_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_285_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_285_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_370 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_383 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_638 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_651 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_732 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_750 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_782 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_308 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_544 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_636 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_705 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1043 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1046 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1052 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1058 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_106 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_286 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_580 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_64 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_788 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_800 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_979 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_187 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_263 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_594 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_711 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_723 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_794 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_896 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_240 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_322 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_519 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_566 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_581 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_763 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_801 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_902 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_914 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_918 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_930 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_942 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_950 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_210 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_292 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_298 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_336 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_399 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_448 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_499 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_575 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_610 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_623 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_631 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_805 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_839 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_860 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_241 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_591 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_614 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_659 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_739 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_815 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_887 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_907 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_919 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_455 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_550 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_568 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_726 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_786 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_826 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_286 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_424 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_496 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_575 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_848 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_854 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_893 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_908 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_932 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_944 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_1093 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_229 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_26 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_280 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_443 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_603 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_680 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_784 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_851 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_857 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_896 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_906 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_971 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_142 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_16 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_413 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_552 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_789 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_804 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_816 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_828 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_84 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_859 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_397 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_678 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_684 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_787 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_873 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_879 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_891 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_899 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_931 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_943 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_955 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_967 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_296 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_39_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_39_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_660 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_39_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_890 ();
 sky130_fd_sc_hd__decap_6 FILLER_39_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_39_920 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_924 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_939 ();
 sky130_fd_sc_hd__fill_1 FILLER_39_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_39_989 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1045 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1056 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1062 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1078 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_130 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_460 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_478 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_688 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_834 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_88 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_246 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_537 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_562 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_654 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_660 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_796 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_40_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_865 ();
 sky130_fd_sc_hd__decap_3 FILLER_40_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_40_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_892 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_904 ();
 sky130_fd_sc_hd__decap_8 FILLER_40_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_40_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_40_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_40_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_10 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_199 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_24 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_63 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_637 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_661 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_41_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_760 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_772 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_779 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_41_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_806 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_846 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_872 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_41_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_41_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_41_910 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_928 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_940 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_41_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_41_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_20 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_298 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_324 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_526 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_732 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_843 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_847 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_42_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_42_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_42_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_42_90 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_42_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_929 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_42_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_42_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_203 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_296 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_308 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_314 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_486 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_496 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_528 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_647 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_725 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_777 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_782 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_799 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_805 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_841 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_863 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_871 ();
 sky130_fd_sc_hd__fill_2 FILLER_43_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_897 ();
 sky130_fd_sc_hd__decap_3 FILLER_43_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_43_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_43_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_43_946 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_43_989 ();
 sky130_fd_sc_hd__decap_8 FILLER_43_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_214 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_224 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_540 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_560 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_44_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_793 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_800 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_44_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_835 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_847 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_44_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_875 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_920 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_44_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_44_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_44_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_44_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_204 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_268 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_410 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_45_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_826 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_832 ();
 sky130_fd_sc_hd__decap_8 FILLER_45_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_853 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_857 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_878 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_890 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_45_945 ();
 sky130_fd_sc_hd__decap_4 FILLER_45_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_45_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_45_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_1093 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_332 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_566 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_635 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_655 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_667 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_822 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_842 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_46_866 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_46_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_904 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_46_916 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_46_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_46_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_46_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_46_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_206 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_47_683 ();
 sky130_fd_sc_hd__decap_3 FILLER_47_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_812 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_864 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_47_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_47_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_911 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_47_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_47_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_47_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_171 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_285 ();
 sky130_fd_sc_hd__decap_3 FILLER_48_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_455 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_462 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_528 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_571 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_606 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_64 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_742 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_820 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_832 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_881 ();
 sky130_fd_sc_hd__decap_8 FILLER_48_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_893 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_911 ();
 sky130_fd_sc_hd__fill_2 FILLER_48_922 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_48_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_48_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_48_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_48_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_140 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_320 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_388 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_527 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_535 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_588 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_49_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_819 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_889 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_912 ();
 sky130_fd_sc_hd__decap_6 FILLER_49_915 ();
 sky130_fd_sc_hd__decap_8 FILLER_49_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_49_949 ();
 sky130_fd_sc_hd__fill_1 FILLER_49_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_49_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_49_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_10 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1049 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1057 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1066 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1080 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1090 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_170 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_272 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_296 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_314 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_576 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_656 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_674 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_684 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_774 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_26 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_381 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_438 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_467 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_572 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_696 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_50_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_776 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_782 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_788 ();
 sky130_fd_sc_hd__decap_3 FILLER_50_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_813 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_819 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_840 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_864 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_894 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_898 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_908 ();
 sky130_fd_sc_hd__decap_4 FILLER_50_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_961 ();
 sky130_fd_sc_hd__decap_6 FILLER_50_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_50_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_50_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_50_997 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_289 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_327 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_35 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_43 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_691 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_774 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_8 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_803 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_809 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_838 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_51_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_856 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_874 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_886 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_894 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_909 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_921 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_51_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_51_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_51_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_51_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_51_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_51_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_618 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_679 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_763 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_784 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_797 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_835 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_841 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_52_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_52_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_902 ();
 sky130_fd_sc_hd__decap_8 FILLER_52_913 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_52_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_52_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_52_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_52_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_254 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_53_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_38 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_409 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_538 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_724 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_745 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_778 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_875 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_882 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_901 ();
 sky130_ef_sc_hd__decap_12 FILLER_53_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_53_925 ();
 sky130_fd_sc_hd__decap_3 FILLER_53_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_53_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_53_98 ();
 sky130_fd_sc_hd__decap_8 FILLER_53_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_117 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_16 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_191 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_414 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_464 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_609 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_761 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_784 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_790 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_798 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_836 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_54_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_854 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_885 ();
 sky130_ef_sc_hd__decap_12 FILLER_54_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_54_942 ();
 sky130_fd_sc_hd__decap_8 FILLER_54_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_54_974 ();
 sky130_fd_sc_hd__decap_3 FILLER_54_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_54_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_241 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_304 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_603 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_55_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_751 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_55_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_823 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_55_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_854 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_906 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_912 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_924 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_55_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_55_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_963 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_55_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_55_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_16 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_355 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_488 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_539 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_791 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_817 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_823 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_840 ();
 sky130_fd_sc_hd__decap_8 FILLER_56_848 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_56_862 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_869 ();
 sky130_fd_sc_hd__decap_3 FILLER_56_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_56_895 ();
 sky130_fd_sc_hd__fill_1 FILLER_56_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_930 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_942 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_954 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_966 ();
 sky130_fd_sc_hd__fill_2 FILLER_56_978 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_56_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1009 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_13 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_149 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_398 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_426 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_438 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_544 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_585 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_57_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_639 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_666 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_72 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_799 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_814 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_841 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_859 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_871 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_894 ();
 sky130_fd_sc_hd__decap_6 FILLER_57_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_911 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_57_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_57_947 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_57_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_975 ();
 sky130_ef_sc_hd__decap_12 FILLER_57_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_57_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1015 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_102 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_138 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_171 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_280 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_416 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_426 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_546 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_63 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_705 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_743 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_780 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_786 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_798 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_810 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_898 ();
 sky130_fd_sc_hd__decap_8 FILLER_58_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_58_91 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_58_932 ();
 sky130_fd_sc_hd__decap_6 FILLER_58_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_941 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_58_965 ();
 sky130_fd_sc_hd__decap_3 FILLER_58_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_58_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_155 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_238 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_298 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_463 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_726 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_752 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_59_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_59_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_831 ();
 sky130_fd_sc_hd__decap_3 FILLER_59_837 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_871 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_59_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_59_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_59_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_59_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1080 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1088 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1098 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1102 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_196 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_310 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_383 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_572 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_753 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_772 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1008 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_20 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_226 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_297 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_379 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_382 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_415 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_550 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_585 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_631 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_731 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_60_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_779 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_785 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_60_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_829 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_910 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_60_932 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_936 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_94 ();
 sky130_fd_sc_hd__decap_8 FILLER_60_960 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_968 ();
 sky130_fd_sc_hd__fill_2 FILLER_60_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_60_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_60_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_37 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_621 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_648 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_756 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_762 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_770 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_61_827 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_885 ();
 sky130_fd_sc_hd__decap_3 FILLER_61_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_61_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_934 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_951 ();
 sky130_fd_sc_hd__decap_6 FILLER_61_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_61_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_61_983 ();
 sky130_fd_sc_hd__decap_8 FILLER_61_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1008 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1020 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_1032 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_1101 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_116 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_124 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_295 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_395 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_467 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_504 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_521 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_58 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_62_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_62_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_848 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_855 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_876 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_62_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_62_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_62_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_974 ();
 sky130_fd_sc_hd__decap_6 FILLER_62_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_62_987 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_266 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_295 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_407 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_479 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_63_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_54 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_723 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_63_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_63_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_63_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_63_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_63_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_63_994 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1010 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1022 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_126 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_20 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_34 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_537 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_625 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_631 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_677 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_720 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_761 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_787 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_64_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_811 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_827 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_848 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_856 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_883 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_64_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_64_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_944 ();
 sky130_fd_sc_hd__decap_8 FILLER_64_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_64_971 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_977 ();
 sky130_fd_sc_hd__decap_3 FILLER_64_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_986 ();
 sky130_ef_sc_hd__decap_12 FILLER_64_998 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_180 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_390 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_466 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_478 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_595 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_700 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_704 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_750 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_758 ();
 sky130_fd_sc_hd__decap_8 FILLER_65_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_811 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_65_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_849 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_894 ();
 sky130_fd_sc_hd__decap_3 FILLER_65_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_926 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_65_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_957 ();
 sky130_fd_sc_hd__fill_1 FILLER_65_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_65_984 ();
 sky130_ef_sc_hd__decap_12 FILLER_65_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1016 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1028 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_12 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_273 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_294 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_361 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_384 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_402 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_452 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_526 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_66_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_619 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_632 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_66_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_750 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_797 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_820 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_834 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_842 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_855 ();
 sky130_fd_sc_hd__decap_6 FILLER_66_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_867 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_66_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_66_938 ();
 sky130_fd_sc_hd__decap_8 FILLER_66_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_66_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_149 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_163 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_219 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_254 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_386 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_419 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_555 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_690 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_721 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_754 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_760 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_67_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_822 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_834 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_864 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_868 ();
 sky130_fd_sc_hd__decap_6 FILLER_67_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_907 ();
 sky130_fd_sc_hd__fill_1 FILLER_67_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_941 ();
 sky130_fd_sc_hd__fill_2 FILLER_67_950 ();
 sky130_fd_sc_hd__decap_3 FILLER_67_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_67_99 ();
 sky130_ef_sc_hd__decap_12 FILLER_67_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1061 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_201 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_230 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_260 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_394 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_436 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_493 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_667 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_68_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_68_787 ();
 sky130_fd_sc_hd__decap_8 FILLER_68_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_8 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_890 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_947 ();
 sky130_fd_sc_hd__decap_6 FILLER_68_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_68_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_68_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_68_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_143 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_201 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_350 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_354 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_408 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_565 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_668 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_695 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_758 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_766 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_772 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_778 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_69_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_69_922 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_928 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_69_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_69_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_962 ();
 sky130_fd_sc_hd__fill_1 FILLER_69_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_972 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_978 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_69_990 ();
 sky130_ef_sc_hd__decap_12 FILLER_69_996 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1083 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1090 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_13 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_271 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_296 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_411 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_509 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_568 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_599 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_611 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_651 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_662 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_731 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_774 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_806 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_156 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_220 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_226 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_24 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_264 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_498 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_510 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_529 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_773 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_779 ();
 sky130_fd_sc_hd__decap_3 FILLER_70_787 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_823 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_829 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_845 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_888 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_912 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_936 ();
 sky130_fd_sc_hd__decap_8 FILLER_70_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_70_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_968 ();
 sky130_fd_sc_hd__decap_6 FILLER_70_974 ();
 sky130_fd_sc_hd__fill_2 FILLER_70_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_70_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_70_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_71_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_200 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_493 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_521 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_617 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_712 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_71_797 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_809 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_835 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_852 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_865 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_941 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_71_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_71_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_71_964 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_71_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_71_999 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_158 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_288 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_338 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_406 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_442 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_450 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_717 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_738 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_744 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_72_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_789 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_72_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_817 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_900 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_916 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_935 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_72_947 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_72_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_72_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_72_991 ();
 sky130_fd_sc_hd__decap_8 FILLER_72_997 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_73_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_158 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_268 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_310 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_332 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_425 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_603 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_622 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_641 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_722 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_73_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_73_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_866 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_73_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_937 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_941 ();
 sky130_fd_sc_hd__decap_6 FILLER_73_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_73_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_73_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_1017 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1023 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_74_1073 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_123 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_389 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_44 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_509 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_530 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_556 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_620 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_697 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_735 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_79 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_799 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_813 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_822 ();
 sky130_fd_sc_hd__fill_1 FILLER_74_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_903 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_929 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_74_963 ();
 sky130_fd_sc_hd__decap_3 FILLER_74_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_74_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_74_985 ();
 sky130_fd_sc_hd__decap_6 FILLER_74_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_75_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_17 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_311 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_323 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_384 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_482 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_75_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_540 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_590 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_633 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_663 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_695 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_751 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_75_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_815 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_825 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_848 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_874 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_890 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_931 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_937 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_946 ();
 sky130_fd_sc_hd__fill_2 FILLER_75_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_966 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_972 ();
 sky130_fd_sc_hd__decap_6 FILLER_75_978 ();
 sky130_fd_sc_hd__fill_1 FILLER_75_984 ();
 sky130_fd_sc_hd__decap_4 FILLER_75_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1026 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1034 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_76_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_194 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_20 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_228 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_34 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_376 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_48 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_527 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_586 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_677 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_723 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_76_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_845 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_893 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_899 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_911 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_923 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_935 ();
 sky130_fd_sc_hd__decap_6 FILLER_76_941 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_947 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_976 ();
 sky130_fd_sc_hd__fill_2 FILLER_76_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_76_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_76_991 ();
 sky130_fd_sc_hd__fill_1 FILLER_76_999 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1006 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_77_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_295 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_316 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_32 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_322 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_446 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_492 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_77_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_567 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_615 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_637 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_664 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_689 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_77_791 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_812 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_77_949 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_95 ();
 sky130_fd_sc_hd__fill_2 FILLER_77_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_77_986 ();
 sky130_fd_sc_hd__decap_6 FILLER_77_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1025 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_103 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_1035 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1053 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_78_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_1089 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_170 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_229 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_330 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_346 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_46 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_506 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_575 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_605 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_631 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_655 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_711 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_717 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_72 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_743 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_776 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_801 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_818 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_847 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_78_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_885 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_944 ();
 sky130_fd_sc_hd__decap_6 FILLER_78_950 ();
 sky130_fd_sc_hd__fill_1 FILLER_78_956 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_78_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_78_985 ();
 sky130_fd_sc_hd__decap_8 FILLER_78_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1036 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1048 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_1060 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_79_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_24 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_30 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_406 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_473 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_522 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_534 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_583 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_604 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_621 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_648 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_782 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_845 ();
 sky130_fd_sc_hd__decap_8 FILLER_79_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_887 ();
 sky130_fd_sc_hd__decap_3 FILLER_79_893 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_912 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_939 ();
 sky130_fd_sc_hd__decap_6 FILLER_79_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_79_951 ();
 sky130_fd_sc_hd__fill_2 FILLER_79_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_968 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_79_995 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1057 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_106 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1077 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1081 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1084 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1095 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_272 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_345 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_351 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_364 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_439 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_581 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_604 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_634 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_659 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_1006 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1030 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_80_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_168 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_17 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_206 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_226 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_263 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_326 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_380 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_431 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_526 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_583 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_612 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_663 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_696 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_719 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_743 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_804 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_810 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_853 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_859 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_865 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_885 ();
 sky130_fd_sc_hd__fill_1 FILLER_80_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_80_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_92 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_947 ();
 sky130_fd_sc_hd__decap_8 FILLER_80_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_80_966 ();
 sky130_fd_sc_hd__decap_3 FILLER_80_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_80_981 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_1005 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1019 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1031 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_81_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_17 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_196 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_232 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_32 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_355 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_358 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_404 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_423 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_430 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_482 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_543 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_649 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_661 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_671 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_719 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_760 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_819 ();
 sky130_fd_sc_hd__fill_1 FILLER_81_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_830 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_836 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_881 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_908 ();
 sky130_fd_sc_hd__decap_8 FILLER_81_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_81_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_81_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_81_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_81_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_82_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_118 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_146 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_22 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_275 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_323 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_34 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_404 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_435 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_472 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_500 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_82_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_562 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_651 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_658 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_664 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_680 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_705 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_781 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_787 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_793 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_811 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_817 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_828 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_834 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_842 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_846 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_856 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_879 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_889 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_902 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_929 ();
 sky130_fd_sc_hd__decap_8 FILLER_82_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_969 ();
 sky130_fd_sc_hd__decap_6 FILLER_82_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_82_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_82_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_985 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_82_997 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1065 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_83_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_173 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_199 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_216 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_243 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_262 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_299 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_34 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_398 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_509 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_592 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_646 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_66 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_695 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_752 ();
 sky130_fd_sc_hd__decap_6 FILLER_83_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_783 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_800 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_806 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_829 ();
 sky130_fd_sc_hd__decap_3 FILLER_83_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_855 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_911 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_922 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_83_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_970 ();
 sky130_fd_sc_hd__decap_4 FILLER_83_976 ();
 sky130_fd_sc_hd__fill_1 FILLER_83_980 ();
 sky130_fd_sc_hd__decap_8 FILLER_83_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1009 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_84_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_145 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_215 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_243 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_249 ();
 sky130_fd_sc_hd__decap_3 FILLER_84_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_276 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_351 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_392 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_428 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_474 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_510 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_522 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_541 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_56 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_564 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_582 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_595 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_616 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_640 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_662 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_676 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_688 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_694 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_780 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_786 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_826 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_839 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_852 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_892 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_899 ();
 sky130_fd_sc_hd__decap_8 FILLER_84_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_906 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_912 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_916 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_84_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_942 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_84_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_979 ();
 sky130_fd_sc_hd__decap_6 FILLER_84_981 ();
 sky130_fd_sc_hd__fill_1 FILLER_84_987 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1077 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_17 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_208 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_258 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_300 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_312 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_341 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_381 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_515 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_547 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_582 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_626 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_85_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_692 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_704 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_715 ();
 sky130_fd_sc_hd__decap_6 FILLER_85_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_795 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_807 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_81 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_818 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_868 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_874 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_880 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_886 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_892 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_919 ();
 sky130_fd_sc_hd__decap_8 FILLER_85_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_85_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_85_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_85_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_85_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_100 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_267 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_304 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_316 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_324 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_327 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_341 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_481 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_58 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_747 ();
 sky130_fd_sc_hd__decap_3 FILLER_86_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_830 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_836 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_842 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_856 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_891 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_903 ();
 sky130_fd_sc_hd__decap_8 FILLER_86_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_920 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_929 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_960 ();
 sky130_fd_sc_hd__decap_4 FILLER_86_966 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_970 ();
 sky130_fd_sc_hd__decap_6 FILLER_86_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_86_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_86_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_86_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_190 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_354 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_381 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_42 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_422 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_457 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_522 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_551 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_557 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_712 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_716 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_87_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_801 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_811 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_827 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_857 ();
 sky130_fd_sc_hd__decap_6 FILLER_87_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_87_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_878 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_884 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_897 ();
 sky130_fd_sc_hd__decap_8 FILLER_87_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_920 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_926 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_938 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_944 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_950 ();
 sky130_fd_sc_hd__fill_2 FILLER_87_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_959 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_87_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_87_995 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_116 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_122 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_228 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_314 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_320 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_349 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_358 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_434 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_531 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_560 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_584 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_661 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_686 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_692 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_706 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_730 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_738 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_747 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_75 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_761 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_794 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_806 ();
 sky130_ef_sc_hd__decap_12 FILLER_88_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_831 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_837 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_849 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_88_855 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_863 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_866 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_892 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_899 ();
 sky130_fd_sc_hd__decap_6 FILLER_88_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_930 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_94 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_942 ();
 sky130_fd_sc_hd__fill_1 FILLER_88_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_967 ();
 sky130_fd_sc_hd__decap_3 FILLER_88_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_88_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_88_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_100 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_1007 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1013 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1025 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1049 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_135 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_183 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_207 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_30 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_310 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_347 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_403 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_435 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_527 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_540 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_89_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_596 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_625 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_638 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_698 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_733 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_774 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_782 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_821 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_845 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_863 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_89_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_887 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_891 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_905 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_916 ();
 sky130_fd_sc_hd__decap_6 FILLER_89_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_927 ();
 sky130_fd_sc_hd__decap_8 FILLER_89_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_89_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_89_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_980 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_89_997 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1029 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_115 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_136 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_230 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_242 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_305 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_322 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_358 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_388 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_394 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_443 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_471 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_606 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_628 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_839 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_881 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_9 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_993 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1000 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1013 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1061 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_1101 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_145 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_231 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_248 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_292 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_303 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_362 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_408 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_427 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_439 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_491 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_523 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_529 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_539 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_547 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_579 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_605 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_62 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_90_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_748 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_767 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_773 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_779 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_791 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_803 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_90_813 ();
 sky130_fd_sc_hd__decap_8 FILLER_90_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_858 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_866 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_869 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_875 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_884 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_896 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_925 ();
 sky130_fd_sc_hd__decap_6 FILLER_90_934 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_959 ();
 sky130_fd_sc_hd__fill_1 FILLER_90_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_90_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_90_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_1004 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_91_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_134 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_160 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_213 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_271 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_28 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_295 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_408 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_466 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_484 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_495 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_524 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_565 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_62 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_623 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_686 ();
 sky130_fd_sc_hd__decap_8 FILLER_91_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_710 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_737 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_773 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_779 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_80 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_802 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_805 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_811 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_839 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_858 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_91_918 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_92 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_937 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_91_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_91_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_969 ();
 sky130_fd_sc_hd__fill_1 FILLER_91_973 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_991 ();
 sky130_fd_sc_hd__decap_4 FILLER_91_998 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1023 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_134 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_192 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_227 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_26 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_294 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_323 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_343 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_356 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_373 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_379 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_385 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_442 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_514 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_520 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_576 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_609 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_667 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_691 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_754 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_768 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_774 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_802 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_810 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_825 ();
 sky130_fd_sc_hd__decap_6 FILLER_92_837 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_864 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_904 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_914 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_940 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_946 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_952 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_959 ();
 sky130_fd_sc_hd__decap_8 FILLER_92_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_92_973 ();
 sky130_fd_sc_hd__decap_3 FILLER_92_977 ();
 sky130_fd_sc_hd__fill_2 FILLER_92_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_92_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_92_999 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_10 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_23 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_245 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_287 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_31 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_390 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_397 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_400 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_467 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_499 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_516 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_542 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_558 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_598 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_607 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_669 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_689 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_694 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_759 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_770 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_776 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_785 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_794 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_809 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_820 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_831 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_850 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_86 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_861 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_872 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_882 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_894 ();
 sky130_fd_sc_hd__decap_8 FILLER_93_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_93_908 ();
 sky130_fd_sc_hd__fill_1 FILLER_93_914 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_917 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_923 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_929 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_943 ();
 sky130_fd_sc_hd__decap_3 FILLER_93_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_93_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_975 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_93_987 ();
 sky130_ef_sc_hd__decap_12 FILLER_93_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_138 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_245 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_25 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_313 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_336 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_362 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_406 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_48 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_582 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_62 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_661 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_667 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_705 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_711 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_72 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_742 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_755 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_803 ();
 sky130_fd_sc_hd__decap_3 FILLER_94_809 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_822 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_833 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_843 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_856 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_869 ();
 sky130_fd_sc_hd__decap_8 FILLER_94_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_906 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_918 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_922 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_925 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_931 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_936 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_943 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_949 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_955 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_961 ();
 sky130_fd_sc_hd__decap_4 FILLER_94_967 ();
 sky130_fd_sc_hd__decap_6 FILLER_94_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_94_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_94_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_985 ();
 sky130_ef_sc_hd__decap_12 FILLER_94_997 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_95_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_140 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_176 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_19 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_222 ();
 sky130_fd_sc_hd__decap_3 FILLER_95_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_334 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_387 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_420 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_423 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_440 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_556 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_590 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_62 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_655 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_659 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_677 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_698 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_726 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_773 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_782 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_785 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_832 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_847 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_859 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_867 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_870 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_876 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_882 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_888 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_907 ();
 sky130_fd_sc_hd__decap_6 FILLER_95_913 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_922 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_935 ();
 sky130_fd_sc_hd__fill_1 FILLER_95_939 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_942 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_948 ();
 sky130_fd_sc_hd__fill_2 FILLER_95_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_957 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_95_993 ();
 sky130_fd_sc_hd__decap_8 FILLER_95_999 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1000 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1012 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1024 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_96_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_1101 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_145 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_148 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_183 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_282 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_306 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_319 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_325 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_328 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_340 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_37 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_400 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_418 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_466 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_533 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_538 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_557 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_628 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_642 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_665 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_68 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_686 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_694 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_730 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_736 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_742 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_748 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_754 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_775 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_799 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_807 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_811 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_821 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_829 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_832 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_838 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_846 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_852 ();
 sky130_fd_sc_hd__decap_6 FILLER_96_858 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_878 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_884 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_890 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_894 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_897 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_901 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_915 ();
 sky130_fd_sc_hd__decap_3 FILLER_96_921 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_925 ();
 sky130_fd_sc_hd__decap_8 FILLER_96_933 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_948 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_954 ();
 sky130_fd_sc_hd__fill_1 FILLER_96_958 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_972 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_96_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_988 ();
 sky130_fd_sc_hd__decap_4 FILLER_96_994 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_1000 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1006 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_1101 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_14 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_187 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_214 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_25 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_348 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_410 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_428 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_443 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_520 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_526 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_565 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_632 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_663 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_682 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_691 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_722 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_775 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_781 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_785 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_792 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_798 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_807 ();
 sky130_ef_sc_hd__decap_12 FILLER_97_813 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_825 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_830 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_834 ();
 sky130_fd_sc_hd__decap_3 FILLER_97_837 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_849 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_857 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_866 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_877 ();
 sky130_fd_sc_hd__decap_8 FILLER_97_883 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_894 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_919 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_932 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_943 ();
 sky130_fd_sc_hd__fill_2 FILLER_97_950 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_953 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_957 ();
 sky130_fd_sc_hd__decap_6 FILLER_97_965 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_979 ();
 sky130_fd_sc_hd__fill_1 FILLER_97_983 ();
 sky130_fd_sc_hd__decap_4 FILLER_97_991 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1003 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1027 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_108 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_1085 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_1091 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_1093 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_114 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_127 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_160 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_184 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_218 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_224 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_285 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_306 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_340 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_344 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_359 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_369 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_372 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_396 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_409 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_485 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_495 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_498 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_504 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_555 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_570 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_58 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_613 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_625 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_675 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_684 ();
 sky130_fd_sc_hd__decap_3 FILLER_98_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_707 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_728 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_734 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_746 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_752 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_761 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_767 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_773 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_777 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_780 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_790 ();
 sky130_ef_sc_hd__decap_12 FILLER_98_796 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_808 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_813 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_817 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_829 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_833 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_844 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_98_856 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_862 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_866 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_873 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_909 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_913 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_922 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_930 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_934 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_943 ();
 sky130_fd_sc_hd__decap_8 FILLER_98_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_954 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_963 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_975 ();
 sky130_fd_sc_hd__fill_1 FILLER_98_979 ();
 sky130_fd_sc_hd__fill_2 FILLER_98_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_98_997 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1002 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_99_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_129 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_203 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_268 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_28 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_36 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_380 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_484 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_496 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_502 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_519 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_543 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_590 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_611 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_654 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_660 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_670 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_688 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_702 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_71 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_718 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_733 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_778 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_789 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_810 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_817 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_828 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_838 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_850 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_860 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_877 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_883 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_895 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_897 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_99_901 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_913 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_924 ();
 sky130_fd_sc_hd__decap_8 FILLER_99_934 ();
 sky130_fd_sc_hd__decap_3 FILLER_99_949 ();
 sky130_fd_sc_hd__fill_2 FILLER_99_953 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_958 ();
 sky130_fd_sc_hd__fill_1 FILLER_99_962 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_969 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_990 ();
 sky130_fd_sc_hd__decap_4 FILLER_99_996 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1033 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1089 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1101 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_117 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_17 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_196 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_230 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_25 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_262 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_269 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_291 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_297 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_355 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_363 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_432 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_438 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_453 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_459 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_465 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_499 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_548 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_578 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_590 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_602 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_794 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_806 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_814 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_818 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_824 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_838 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_855 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_867 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_879 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_887 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_977 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_989 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_314 ();
 sky130_fd_sc_hd__decap_3 PHY_315 ();
 sky130_fd_sc_hd__decap_3 PHY_316 ();
 sky130_fd_sc_hd__decap_3 PHY_317 ();
 sky130_fd_sc_hd__decap_3 PHY_318 ();
 sky130_fd_sc_hd__decap_3 PHY_319 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_320 ();
 sky130_fd_sc_hd__decap_3 PHY_321 ();
 sky130_fd_sc_hd__decap_3 PHY_322 ();
 sky130_fd_sc_hd__decap_3 PHY_323 ();
 sky130_fd_sc_hd__decap_3 PHY_324 ();
 sky130_fd_sc_hd__decap_3 PHY_325 ();
 sky130_fd_sc_hd__decap_3 PHY_326 ();
 sky130_fd_sc_hd__decap_3 PHY_327 ();
 sky130_fd_sc_hd__decap_3 PHY_328 ();
 sky130_fd_sc_hd__decap_3 PHY_329 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_330 ();
 sky130_fd_sc_hd__decap_3 PHY_331 ();
 sky130_fd_sc_hd__decap_3 PHY_332 ();
 sky130_fd_sc_hd__decap_3 PHY_333 ();
 sky130_fd_sc_hd__decap_3 PHY_334 ();
 sky130_fd_sc_hd__decap_3 PHY_335 ();
 sky130_fd_sc_hd__decap_3 PHY_336 ();
 sky130_fd_sc_hd__decap_3 PHY_337 ();
 sky130_fd_sc_hd__decap_3 PHY_338 ();
 sky130_fd_sc_hd__decap_3 PHY_339 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_340 ();
 sky130_fd_sc_hd__decap_3 PHY_341 ();
 sky130_fd_sc_hd__decap_3 PHY_342 ();
 sky130_fd_sc_hd__decap_3 PHY_343 ();
 sky130_fd_sc_hd__decap_3 PHY_344 ();
 sky130_fd_sc_hd__decap_3 PHY_345 ();
 sky130_fd_sc_hd__decap_3 PHY_346 ();
 sky130_fd_sc_hd__decap_3 PHY_347 ();
 sky130_fd_sc_hd__decap_3 PHY_348 ();
 sky130_fd_sc_hd__decap_3 PHY_349 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_350 ();
 sky130_fd_sc_hd__decap_3 PHY_351 ();
 sky130_fd_sc_hd__decap_3 PHY_352 ();
 sky130_fd_sc_hd__decap_3 PHY_353 ();
 sky130_fd_sc_hd__decap_3 PHY_354 ();
 sky130_fd_sc_hd__decap_3 PHY_355 ();
 sky130_fd_sc_hd__decap_3 PHY_356 ();
 sky130_fd_sc_hd__decap_3 PHY_357 ();
 sky130_fd_sc_hd__decap_3 PHY_358 ();
 sky130_fd_sc_hd__decap_3 PHY_359 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_360 ();
 sky130_fd_sc_hd__decap_3 PHY_361 ();
 sky130_fd_sc_hd__decap_3 PHY_362 ();
 sky130_fd_sc_hd__decap_3 PHY_363 ();
 sky130_fd_sc_hd__decap_3 PHY_364 ();
 sky130_fd_sc_hd__decap_3 PHY_365 ();
 sky130_fd_sc_hd__decap_3 PHY_366 ();
 sky130_fd_sc_hd__decap_3 PHY_367 ();
 sky130_fd_sc_hd__decap_3 PHY_368 ();
 sky130_fd_sc_hd__decap_3 PHY_369 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_370 ();
 sky130_fd_sc_hd__decap_3 PHY_371 ();
 sky130_fd_sc_hd__decap_3 PHY_372 ();
 sky130_fd_sc_hd__decap_3 PHY_373 ();
 sky130_fd_sc_hd__decap_3 PHY_374 ();
 sky130_fd_sc_hd__decap_3 PHY_375 ();
 sky130_fd_sc_hd__decap_3 PHY_376 ();
 sky130_fd_sc_hd__decap_3 PHY_377 ();
 sky130_fd_sc_hd__decap_3 PHY_378 ();
 sky130_fd_sc_hd__decap_3 PHY_379 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_380 ();
 sky130_fd_sc_hd__decap_3 PHY_381 ();
 sky130_fd_sc_hd__decap_3 PHY_382 ();
 sky130_fd_sc_hd__decap_3 PHY_383 ();
 sky130_fd_sc_hd__decap_3 PHY_384 ();
 sky130_fd_sc_hd__decap_3 PHY_385 ();
 sky130_fd_sc_hd__decap_3 PHY_386 ();
 sky130_fd_sc_hd__decap_3 PHY_387 ();
 sky130_fd_sc_hd__decap_3 PHY_388 ();
 sky130_fd_sc_hd__decap_3 PHY_389 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_390 ();
 sky130_fd_sc_hd__decap_3 PHY_391 ();
 sky130_fd_sc_hd__decap_3 PHY_392 ();
 sky130_fd_sc_hd__decap_3 PHY_393 ();
 sky130_fd_sc_hd__decap_3 PHY_394 ();
 sky130_fd_sc_hd__decap_3 PHY_395 ();
 sky130_fd_sc_hd__decap_3 PHY_396 ();
 sky130_fd_sc_hd__decap_3 PHY_397 ();
 sky130_fd_sc_hd__decap_3 PHY_398 ();
 sky130_fd_sc_hd__decap_3 PHY_399 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_400 ();
 sky130_fd_sc_hd__decap_3 PHY_401 ();
 sky130_fd_sc_hd__decap_3 PHY_402 ();
 sky130_fd_sc_hd__decap_3 PHY_403 ();
 sky130_fd_sc_hd__decap_3 PHY_404 ();
 sky130_fd_sc_hd__decap_3 PHY_405 ();
 sky130_fd_sc_hd__decap_3 PHY_406 ();
 sky130_fd_sc_hd__decap_3 PHY_407 ();
 sky130_fd_sc_hd__decap_3 PHY_408 ();
 sky130_fd_sc_hd__decap_3 PHY_409 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_410 ();
 sky130_fd_sc_hd__decap_3 PHY_411 ();
 sky130_fd_sc_hd__decap_3 PHY_412 ();
 sky130_fd_sc_hd__decap_3 PHY_413 ();
 sky130_fd_sc_hd__decap_3 PHY_414 ();
 sky130_fd_sc_hd__decap_3 PHY_415 ();
 sky130_fd_sc_hd__decap_3 PHY_416 ();
 sky130_fd_sc_hd__decap_3 PHY_417 ();
 sky130_fd_sc_hd__decap_3 PHY_418 ();
 sky130_fd_sc_hd__decap_3 PHY_419 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_420 ();
 sky130_fd_sc_hd__decap_3 PHY_421 ();
 sky130_fd_sc_hd__decap_3 PHY_422 ();
 sky130_fd_sc_hd__decap_3 PHY_423 ();
 sky130_fd_sc_hd__decap_3 PHY_424 ();
 sky130_fd_sc_hd__decap_3 PHY_425 ();
 sky130_fd_sc_hd__decap_3 PHY_426 ();
 sky130_fd_sc_hd__decap_3 PHY_427 ();
 sky130_fd_sc_hd__decap_3 PHY_428 ();
 sky130_fd_sc_hd__decap_3 PHY_429 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_430 ();
 sky130_fd_sc_hd__decap_3 PHY_431 ();
 sky130_fd_sc_hd__decap_3 PHY_432 ();
 sky130_fd_sc_hd__decap_3 PHY_433 ();
 sky130_fd_sc_hd__decap_3 PHY_434 ();
 sky130_fd_sc_hd__decap_3 PHY_435 ();
 sky130_fd_sc_hd__decap_3 PHY_436 ();
 sky130_fd_sc_hd__decap_3 PHY_437 ();
 sky130_fd_sc_hd__decap_3 PHY_438 ();
 sky130_fd_sc_hd__decap_3 PHY_439 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_440 ();
 sky130_fd_sc_hd__decap_3 PHY_441 ();
 sky130_fd_sc_hd__decap_3 PHY_442 ();
 sky130_fd_sc_hd__decap_3 PHY_443 ();
 sky130_fd_sc_hd__decap_3 PHY_444 ();
 sky130_fd_sc_hd__decap_3 PHY_445 ();
 sky130_fd_sc_hd__decap_3 PHY_446 ();
 sky130_fd_sc_hd__decap_3 PHY_447 ();
 sky130_fd_sc_hd__decap_3 PHY_448 ();
 sky130_fd_sc_hd__decap_3 PHY_449 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_450 ();
 sky130_fd_sc_hd__decap_3 PHY_451 ();
 sky130_fd_sc_hd__decap_3 PHY_452 ();
 sky130_fd_sc_hd__decap_3 PHY_453 ();
 sky130_fd_sc_hd__decap_3 PHY_454 ();
 sky130_fd_sc_hd__decap_3 PHY_455 ();
 sky130_fd_sc_hd__decap_3 PHY_456 ();
 sky130_fd_sc_hd__decap_3 PHY_457 ();
 sky130_fd_sc_hd__decap_3 PHY_458 ();
 sky130_fd_sc_hd__decap_3 PHY_459 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_460 ();
 sky130_fd_sc_hd__decap_3 PHY_461 ();
 sky130_fd_sc_hd__decap_3 PHY_462 ();
 sky130_fd_sc_hd__decap_3 PHY_463 ();
 sky130_fd_sc_hd__decap_3 PHY_464 ();
 sky130_fd_sc_hd__decap_3 PHY_465 ();
 sky130_fd_sc_hd__decap_3 PHY_466 ();
 sky130_fd_sc_hd__decap_3 PHY_467 ();
 sky130_fd_sc_hd__decap_3 PHY_468 ();
 sky130_fd_sc_hd__decap_3 PHY_469 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_470 ();
 sky130_fd_sc_hd__decap_3 PHY_471 ();
 sky130_fd_sc_hd__decap_3 PHY_472 ();
 sky130_fd_sc_hd__decap_3 PHY_473 ();
 sky130_fd_sc_hd__decap_3 PHY_474 ();
 sky130_fd_sc_hd__decap_3 PHY_475 ();
 sky130_fd_sc_hd__decap_3 PHY_476 ();
 sky130_fd_sc_hd__decap_3 PHY_477 ();
 sky130_fd_sc_hd__decap_3 PHY_478 ();
 sky130_fd_sc_hd__decap_3 PHY_479 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_480 ();
 sky130_fd_sc_hd__decap_3 PHY_481 ();
 sky130_fd_sc_hd__decap_3 PHY_482 ();
 sky130_fd_sc_hd__decap_3 PHY_483 ();
 sky130_fd_sc_hd__decap_3 PHY_484 ();
 sky130_fd_sc_hd__decap_3 PHY_485 ();
 sky130_fd_sc_hd__decap_3 PHY_486 ();
 sky130_fd_sc_hd__decap_3 PHY_487 ();
 sky130_fd_sc_hd__decap_3 PHY_488 ();
 sky130_fd_sc_hd__decap_3 PHY_489 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_490 ();
 sky130_fd_sc_hd__decap_3 PHY_491 ();
 sky130_fd_sc_hd__decap_3 PHY_492 ();
 sky130_fd_sc_hd__decap_3 PHY_493 ();
 sky130_fd_sc_hd__decap_3 PHY_494 ();
 sky130_fd_sc_hd__decap_3 PHY_495 ();
 sky130_fd_sc_hd__decap_3 PHY_496 ();
 sky130_fd_sc_hd__decap_3 PHY_497 ();
 sky130_fd_sc_hd__decap_3 PHY_498 ();
 sky130_fd_sc_hd__decap_3 PHY_499 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_500 ();
 sky130_fd_sc_hd__decap_3 PHY_501 ();
 sky130_fd_sc_hd__decap_3 PHY_502 ();
 sky130_fd_sc_hd__decap_3 PHY_503 ();
 sky130_fd_sc_hd__decap_3 PHY_504 ();
 sky130_fd_sc_hd__decap_3 PHY_505 ();
 sky130_fd_sc_hd__decap_3 PHY_506 ();
 sky130_fd_sc_hd__decap_3 PHY_507 ();
 sky130_fd_sc_hd__decap_3 PHY_508 ();
 sky130_fd_sc_hd__decap_3 PHY_509 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_510 ();
 sky130_fd_sc_hd__decap_3 PHY_511 ();
 sky130_fd_sc_hd__decap_3 PHY_512 ();
 sky130_fd_sc_hd__decap_3 PHY_513 ();
 sky130_fd_sc_hd__decap_3 PHY_514 ();
 sky130_fd_sc_hd__decap_3 PHY_515 ();
 sky130_fd_sc_hd__decap_3 PHY_516 ();
 sky130_fd_sc_hd__decap_3 PHY_517 ();
 sky130_fd_sc_hd__decap_3 PHY_518 ();
 sky130_fd_sc_hd__decap_3 PHY_519 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_520 ();
 sky130_fd_sc_hd__decap_3 PHY_521 ();
 sky130_fd_sc_hd__decap_3 PHY_522 ();
 sky130_fd_sc_hd__decap_3 PHY_523 ();
 sky130_fd_sc_hd__decap_3 PHY_524 ();
 sky130_fd_sc_hd__decap_3 PHY_525 ();
 sky130_fd_sc_hd__decap_3 PHY_526 ();
 sky130_fd_sc_hd__decap_3 PHY_527 ();
 sky130_fd_sc_hd__decap_3 PHY_528 ();
 sky130_fd_sc_hd__decap_3 PHY_529 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_530 ();
 sky130_fd_sc_hd__decap_3 PHY_531 ();
 sky130_fd_sc_hd__decap_3 PHY_532 ();
 sky130_fd_sc_hd__decap_3 PHY_533 ();
 sky130_fd_sc_hd__decap_3 PHY_534 ();
 sky130_fd_sc_hd__decap_3 PHY_535 ();
 sky130_fd_sc_hd__decap_3 PHY_536 ();
 sky130_fd_sc_hd__decap_3 PHY_537 ();
 sky130_fd_sc_hd__decap_3 PHY_538 ();
 sky130_fd_sc_hd__decap_3 PHY_539 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_540 ();
 sky130_fd_sc_hd__decap_3 PHY_541 ();
 sky130_fd_sc_hd__decap_3 PHY_542 ();
 sky130_fd_sc_hd__decap_3 PHY_543 ();
 sky130_fd_sc_hd__decap_3 PHY_544 ();
 sky130_fd_sc_hd__decap_3 PHY_545 ();
 sky130_fd_sc_hd__decap_3 PHY_546 ();
 sky130_fd_sc_hd__decap_3 PHY_547 ();
 sky130_fd_sc_hd__decap_3 PHY_548 ();
 sky130_fd_sc_hd__decap_3 PHY_549 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_550 ();
 sky130_fd_sc_hd__decap_3 PHY_551 ();
 sky130_fd_sc_hd__decap_3 PHY_552 ();
 sky130_fd_sc_hd__decap_3 PHY_553 ();
 sky130_fd_sc_hd__decap_3 PHY_554 ();
 sky130_fd_sc_hd__decap_3 PHY_555 ();
 sky130_fd_sc_hd__decap_3 PHY_556 ();
 sky130_fd_sc_hd__decap_3 PHY_557 ();
 sky130_fd_sc_hd__decap_3 PHY_558 ();
 sky130_fd_sc_hd__decap_3 PHY_559 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_560 ();
 sky130_fd_sc_hd__decap_3 PHY_561 ();
 sky130_fd_sc_hd__decap_3 PHY_562 ();
 sky130_fd_sc_hd__decap_3 PHY_563 ();
 sky130_fd_sc_hd__decap_3 PHY_564 ();
 sky130_fd_sc_hd__decap_3 PHY_565 ();
 sky130_fd_sc_hd__decap_3 PHY_566 ();
 sky130_fd_sc_hd__decap_3 PHY_567 ();
 sky130_fd_sc_hd__decap_3 PHY_568 ();
 sky130_fd_sc_hd__decap_3 PHY_569 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_570 ();
 sky130_fd_sc_hd__decap_3 PHY_571 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_3999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_4999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_5999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_6187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _04688_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.wr_ptr ),
    .Y(_04343_));
 sky130_fd_sc_hd__inv_2 _04689_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.wr_ptr ),
    .Y(_04345_));
 sky130_fd_sc_hd__clkinv_2 _04690_ (.A(net1084),
    .Y(_04346_));
 sky130_fd_sc_hd__inv_2 _04691_ (.A(net130),
    .Y(_00776_));
 sky130_fd_sc_hd__inv_2 _04692_ (.A(net1348),
    .Y(_00777_));
 sky130_fd_sc_hd__inv_2 _04693_ (.A(net1368),
    .Y(_00778_));
 sky130_fd_sc_hd__inv_2 _04694_ (.A(net1345),
    .Y(_00779_));
 sky130_fd_sc_hd__inv_2 _04695_ (.A(\u_gpio.u_bit[10].u_dglitch.gpio_reg ),
    .Y(_00780_));
 sky130_fd_sc_hd__inv_2 _04696_ (.A(\u_gpio.u_bit[11].u_dglitch.gpio_reg ),
    .Y(_00781_));
 sky130_fd_sc_hd__inv_2 _04697_ (.A(\u_gpio.u_bit[12].u_dglitch.gpio_reg ),
    .Y(_00782_));
 sky130_fd_sc_hd__inv_2 _04698_ (.A(\u_gpio.u_bit[13].u_dglitch.gpio_reg ),
    .Y(_00783_));
 sky130_fd_sc_hd__inv_2 _04699_ (.A(\u_gpio.u_bit[14].u_dglitch.gpio_reg ),
    .Y(_00784_));
 sky130_fd_sc_hd__inv_2 _04700_ (.A(\u_gpio.u_bit[15].u_dglitch.gpio_reg ),
    .Y(_00785_));
 sky130_fd_sc_hd__inv_2 _04701_ (.A(\u_gpio.u_bit[16].u_dglitch.gpio_reg ),
    .Y(_00786_));
 sky130_fd_sc_hd__inv_2 _04702_ (.A(\u_gpio.u_bit[17].u_dglitch.gpio_reg ),
    .Y(_00787_));
 sky130_fd_sc_hd__inv_2 _04703_ (.A(\u_gpio.u_bit[18].u_dglitch.gpio_reg ),
    .Y(_00788_));
 sky130_fd_sc_hd__inv_2 _04704_ (.A(\u_gpio.u_bit[20].u_dglitch.gpio_reg ),
    .Y(_00789_));
 sky130_fd_sc_hd__inv_2 _04705_ (.A(\u_gpio.u_bit[21].u_dglitch.gpio_reg ),
    .Y(_00790_));
 sky130_fd_sc_hd__inv_2 _04706_ (.A(\u_gpio.u_bit[22].u_dglitch.gpio_reg ),
    .Y(_00791_));
 sky130_fd_sc_hd__inv_2 _04707_ (.A(\u_gpio.u_bit[8].u_dglitch.gpio_reg ),
    .Y(_00792_));
 sky130_fd_sc_hd__inv_2 _04708_ (.A(\u_gpio.u_bit[9].u_dglitch.gpio_reg ),
    .Y(_00793_));
 sky130_fd_sc_hd__clkinv_2 _04709_ (.A(\u_glbl_reg.u_dbgclk.high_count[0] ),
    .Y(_00039_));
 sky130_fd_sc_hd__inv_2 _04710_ (.A(net1343),
    .Y(_00794_));
 sky130_fd_sc_hd__inv_2 _04711_ (.A(net774),
    .Y(_00795_));
 sky130_fd_sc_hd__inv_2 _04712_ (.A(net1055),
    .Y(_00796_));
 sky130_fd_sc_hd__inv_2 _04713_ (.A(\u_ws281x.cfg_clk_period[0] ),
    .Y(_00797_));
 sky130_fd_sc_hd__clkinv_2 _04714_ (.A(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .Y(_00798_));
 sky130_fd_sc_hd__inv_2 _04715_ (.A(\u_ws281x.cfg_clk_period[1] ),
    .Y(_00799_));
 sky130_fd_sc_hd__inv_2 _04716_ (.A(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .Y(_00800_));
 sky130_fd_sc_hd__inv_2 _04717_ (.A(\u_ws281x.cfg_clk_period[2] ),
    .Y(_00801_));
 sky130_fd_sc_hd__clkinv_2 _04718_ (.A(\u_ws281x.u_txd_0.clk_cnt[2] ),
    .Y(_00802_));
 sky130_fd_sc_hd__inv_2 _04719_ (.A(\u_ws281x.cfg_clk_period[3] ),
    .Y(_00803_));
 sky130_fd_sc_hd__clkinv_2 _04720_ (.A(\u_ws281x.u_txd_0.clk_cnt[3] ),
    .Y(_00804_));
 sky130_fd_sc_hd__clkinv_2 _04721_ (.A(\u_ws281x.u_txd_0.clk_cnt[4] ),
    .Y(_00805_));
 sky130_fd_sc_hd__inv_2 _04722_ (.A(\u_ws281x.cfg_clk_period[5] ),
    .Y(_00806_));
 sky130_fd_sc_hd__inv_2 _04723_ (.A(\u_ws281x.u_txd_0.clk_cnt[5] ),
    .Y(_00807_));
 sky130_fd_sc_hd__clkinv_2 _04724_ (.A(\u_ws281x.u_txd_0.clk_cnt[6] ),
    .Y(_00808_));
 sky130_fd_sc_hd__inv_2 _04725_ (.A(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .Y(_00809_));
 sky130_fd_sc_hd__inv_2 _04726_ (.A(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .Y(_00810_));
 sky130_fd_sc_hd__inv_2 _04727_ (.A(\u_ws281x.cfg_clk_period[9] ),
    .Y(_00811_));
 sky130_fd_sc_hd__inv_2 _04728_ (.A(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .Y(_00812_));
 sky130_fd_sc_hd__inv_2 _04729_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .Y(_00813_));
 sky130_fd_sc_hd__inv_2 _04730_ (.A(\u_ws281x.cfg_reset_period[1] ),
    .Y(_00814_));
 sky130_fd_sc_hd__inv_2 _04731_ (.A(\u_ws281x.cfg_reset_period[3] ),
    .Y(_00815_));
 sky130_fd_sc_hd__inv_2 _04732_ (.A(\u_ws281x.cfg_reset_period[5] ),
    .Y(_00816_));
 sky130_fd_sc_hd__inv_2 _04733_ (.A(\u_ws281x.cfg_reset_period[6] ),
    .Y(_00817_));
 sky130_fd_sc_hd__inv_2 _04734_ (.A(\u_ws281x.cfg_reset_period[7] ),
    .Y(_00818_));
 sky130_fd_sc_hd__inv_2 _04735_ (.A(\u_ws281x.cfg_reset_period[8] ),
    .Y(_00819_));
 sky130_fd_sc_hd__inv_2 _04736_ (.A(\u_ws281x.cfg_reset_period[9] ),
    .Y(_00820_));
 sky130_fd_sc_hd__inv_2 _04737_ (.A(\u_ws281x.cfg_reset_period[11] ),
    .Y(_00821_));
 sky130_fd_sc_hd__inv_2 _04738_ (.A(\u_ws281x.cfg_reset_period[12] ),
    .Y(_00822_));
 sky130_fd_sc_hd__inv_2 _04739_ (.A(\u_ws281x.cfg_reset_period[13] ),
    .Y(_00823_));
 sky130_fd_sc_hd__inv_2 _04740_ (.A(\u_ws281x.cfg_reset_period[15] ),
    .Y(_00824_));
 sky130_fd_sc_hd__inv_2 _04741_ (.A(net2342),
    .Y(_00825_));
 sky130_fd_sc_hd__clkinv_2 _04742_ (.A(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .Y(_00826_));
 sky130_fd_sc_hd__inv_2 _04743_ (.A(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .Y(_00827_));
 sky130_fd_sc_hd__clkinv_2 _04744_ (.A(\u_ws281x.u_txd_1.clk_cnt[2] ),
    .Y(_00828_));
 sky130_fd_sc_hd__clkinv_2 _04745_ (.A(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .Y(_00829_));
 sky130_fd_sc_hd__clkinv_2 _04746_ (.A(\u_ws281x.u_txd_1.clk_cnt[4] ),
    .Y(_00830_));
 sky130_fd_sc_hd__inv_2 _04747_ (.A(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .Y(_00831_));
 sky130_fd_sc_hd__clkinv_2 _04748_ (.A(\u_ws281x.u_txd_1.clk_cnt[6] ),
    .Y(_00832_));
 sky130_fd_sc_hd__inv_2 _04749_ (.A(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .Y(_00833_));
 sky130_fd_sc_hd__clkinv_2 _04750_ (.A(\u_ws281x.u_txd_1.clk_cnt[8] ),
    .Y(_00834_));
 sky130_fd_sc_hd__inv_2 _04751_ (.A(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .Y(_00835_));
 sky130_fd_sc_hd__inv_2 _04752_ (.A(\u_ws281x.u_txd_1.clk_cnt[11] ),
    .Y(_00836_));
 sky130_fd_sc_hd__inv_2 _04753_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .Y(_00837_));
 sky130_fd_sc_hd__inv_2 _04754_ (.A(\u_ws281x.port1_enb ),
    .Y(_00838_));
 sky130_fd_sc_hd__inv_2 _04755_ (.A(net2348),
    .Y(_00839_));
 sky130_fd_sc_hd__clkinv_2 _04756_ (.A(\u_timer.u_timer_2.timer_counter[0] ),
    .Y(_00840_));
 sky130_fd_sc_hd__inv_2 _04757_ (.A(\u_timer.u_timer_2.timer_hit_s1 ),
    .Y(_00841_));
 sky130_fd_sc_hd__inv_2 _04758_ (.A(\u_timer.cfg_timer2[16] ),
    .Y(_00842_));
 sky130_fd_sc_hd__clkinv_2 _04759_ (.A(\u_timer.u_timer_1.timer_counter[0] ),
    .Y(_00843_));
 sky130_fd_sc_hd__inv_2 _04760_ (.A(\u_timer.u_timer_1.timer_hit_s1 ),
    .Y(_00844_));
 sky130_fd_sc_hd__inv_2 _04761_ (.A(\u_timer.cfg_timer1[16] ),
    .Y(_00845_));
 sky130_fd_sc_hd__clkinv_2 _04762_ (.A(\u_timer.u_timer_0.timer_counter[0] ),
    .Y(_00846_));
 sky130_fd_sc_hd__inv_2 _04763_ (.A(\u_timer.u_timer_0.timer_hit_s1 ),
    .Y(_00847_));
 sky130_fd_sc_hd__inv_2 _04764_ (.A(\u_timer.cfg_timer0[16] ),
    .Y(_00848_));
 sky130_fd_sc_hd__inv_2 _04765_ (.A(\u_ws281x.port1_rd ),
    .Y(_00849_));
 sky130_fd_sc_hd__inv_2 _04766_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.full ),
    .Y(_00850_));
 sky130_fd_sc_hd__inv_2 _04767_ (.A(\u_ws281x.port0_rd ),
    .Y(_00851_));
 sky130_fd_sc_hd__clkinv_2 _04768_ (.A(net1080),
    .Y(_04344_));
 sky130_fd_sc_hd__inv_2 _04769_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.full ),
    .Y(_00852_));
 sky130_fd_sc_hd__inv_2 _04770_ (.A(\u_ws281x.cfg_th0_period[9] ),
    .Y(_00853_));
 sky130_fd_sc_hd__inv_2 _04771_ (.A(\u_ws281x.cfg_th1_period[3] ),
    .Y(_00854_));
 sky130_fd_sc_hd__inv_2 _04772_ (.A(\u_ws281x.cfg_th1_period[7] ),
    .Y(_00855_));
 sky130_fd_sc_hd__inv_2 _04773_ (.A(\u_timer.u_pulse_1ms.cnt[9] ),
    .Y(_00856_));
 sky130_fd_sc_hd__inv_2 _04774_ (.A(\u_timer.u_pulse_1s.cnt[9] ),
    .Y(_00857_));
 sky130_fd_sc_hd__inv_2 _04775_ (.A(net1076),
    .Y(_00858_));
 sky130_fd_sc_hd__clkinv_2 _04776_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .Y(_00859_));
 sky130_fd_sc_hd__inv_2 _04777_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .Y(_00860_));
 sky130_fd_sc_hd__clkinv_2 _04778_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .Y(_00861_));
 sky130_fd_sc_hd__clkinv_2 _04779_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .Y(_00862_));
 sky130_fd_sc_hd__clkinv_2 _04780_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .Y(_00863_));
 sky130_fd_sc_hd__inv_2 _04781_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .Y(_00864_));
 sky130_fd_sc_hd__inv_2 _04782_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ),
    .Y(_00865_));
 sky130_fd_sc_hd__inv_2 _04783_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .Y(_00866_));
 sky130_fd_sc_hd__inv_2 _04784_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ),
    .Y(_00867_));
 sky130_fd_sc_hd__inv_2 _04785_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ),
    .Y(_00868_));
 sky130_fd_sc_hd__inv_2 _04786_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .Y(_00869_));
 sky130_fd_sc_hd__inv_2 _04787_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ),
    .Y(_00870_));
 sky130_fd_sc_hd__inv_2 _04788_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ),
    .Y(_00871_));
 sky130_fd_sc_hd__inv_2 _04789_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .Y(_00872_));
 sky130_fd_sc_hd__clkinv_2 _04790_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .Y(_00873_));
 sky130_fd_sc_hd__inv_2 _04791_ (.A(\u_pwm.u_pwm_0.cfg_pwm_period[3] ),
    .Y(_00874_));
 sky130_fd_sc_hd__inv_2 _04792_ (.A(\u_pwm.u_pwm_0.cfg_pwm_period[11] ),
    .Y(_00875_));
 sky130_fd_sc_hd__inv_2 _04793_ (.A(\u_pwm.u_pwm_0.cfg_pwm_period[12] ),
    .Y(_00876_));
 sky130_fd_sc_hd__inv_2 _04794_ (.A(\u_pwm.u_pwm_0.cfg_pwm_period[13] ),
    .Y(_00877_));
 sky130_fd_sc_hd__inv_2 _04795_ (.A(net1075),
    .Y(_00878_));
 sky130_fd_sc_hd__clkinv_2 _04796_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .Y(_00879_));
 sky130_fd_sc_hd__clkinv_2 _04797_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .Y(_00880_));
 sky130_fd_sc_hd__clkinv_2 _04798_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .Y(_00881_));
 sky130_fd_sc_hd__clkinv_2 _04799_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .Y(_00882_));
 sky130_fd_sc_hd__inv_2 _04800_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .Y(_00883_));
 sky130_fd_sc_hd__clkinv_2 _04801_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .Y(_00884_));
 sky130_fd_sc_hd__clkinv_4 _04802_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ),
    .Y(_00885_));
 sky130_fd_sc_hd__inv_2 _04803_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ),
    .Y(_00886_));
 sky130_fd_sc_hd__inv_2 _04804_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ),
    .Y(_00887_));
 sky130_fd_sc_hd__inv_2 _04805_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[5] ),
    .Y(_00888_));
 sky130_fd_sc_hd__inv_2 _04806_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .Y(_00889_));
 sky130_fd_sc_hd__clkinv_2 _04807_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .Y(_00890_));
 sky130_fd_sc_hd__inv_2 _04808_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .Y(_00891_));
 sky130_fd_sc_hd__clkinv_2 _04809_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .Y(_00892_));
 sky130_fd_sc_hd__clkinv_2 _04810_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .Y(_00893_));
 sky130_fd_sc_hd__inv_2 _04811_ (.A(\u_pwm.u_pwm_1.cfg_pwm_period[0] ),
    .Y(_00894_));
 sky130_fd_sc_hd__inv_2 _04812_ (.A(\u_pwm.u_pwm_1.cfg_pwm_period[1] ),
    .Y(_00895_));
 sky130_fd_sc_hd__inv_2 _04813_ (.A(\u_pwm.u_pwm_1.cfg_pwm_period[3] ),
    .Y(_00896_));
 sky130_fd_sc_hd__inv_2 _04814_ (.A(\u_pwm.u_pwm_1.cfg_pwm_period[11] ),
    .Y(_00897_));
 sky130_fd_sc_hd__inv_2 _04815_ (.A(net1071),
    .Y(_00898_));
 sky130_fd_sc_hd__clkinv_2 _04816_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[14] ),
    .Y(_00899_));
 sky130_fd_sc_hd__clkinv_2 _04817_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .Y(_00900_));
 sky130_fd_sc_hd__clkinv_2 _04818_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .Y(_00901_));
 sky130_fd_sc_hd__clkinv_2 _04819_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .Y(_00902_));
 sky130_fd_sc_hd__inv_2 _04820_ (.A(net1073),
    .Y(_00903_));
 sky130_fd_sc_hd__inv_2 _04821_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .Y(_00904_));
 sky130_fd_sc_hd__clkinv_2 _04822_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .Y(_00905_));
 sky130_fd_sc_hd__inv_2 _04823_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .Y(_00906_));
 sky130_fd_sc_hd__clkinv_2 _04824_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .Y(_00907_));
 sky130_fd_sc_hd__inv_2 _04825_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ),
    .Y(_00908_));
 sky130_fd_sc_hd__clkinv_2 _04826_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .Y(_00909_));
 sky130_fd_sc_hd__inv_2 _04827_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ),
    .Y(_00910_));
 sky130_fd_sc_hd__inv_2 _04828_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ),
    .Y(_00911_));
 sky130_fd_sc_hd__clkinv_2 _04829_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .Y(_00912_));
 sky130_fd_sc_hd__clkinv_2 _04830_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ),
    .Y(_00913_));
 sky130_fd_sc_hd__inv_2 _04831_ (.A(\u_pwm.u_pwm_2.cfg_pwm_period[4] ),
    .Y(_00914_));
 sky130_fd_sc_hd__inv_2 _04832_ (.A(\u_pwm.u_pwm_2.cfg_pwm_period[11] ),
    .Y(_00915_));
 sky130_fd_sc_hd__inv_2 _04833_ (.A(\u_pwm.u_pwm_2.cfg_pwm_period[12] ),
    .Y(_00916_));
 sky130_fd_sc_hd__inv_2 _04834_ (.A(\u_pwm.u_pwm_2.cfg_pwm_period[13] ),
    .Y(_00917_));
 sky130_fd_sc_hd__inv_2 _04835_ (.A(\u_pwm.u_pwm_0.cfg_pwm_scale[2] ),
    .Y(_00918_));
 sky130_fd_sc_hd__inv_2 _04836_ (.A(\u_pwm.u_pwm_0.cfg_pwm_scale[0] ),
    .Y(_00919_));
 sky130_fd_sc_hd__inv_2 _04837_ (.A(\u_pwm.u_pwm_0.cfg_pwm_scale[1] ),
    .Y(_00920_));
 sky130_fd_sc_hd__inv_2 _04838_ (.A(\u_pwm.u_pwm_1.cfg_pwm_scale[2] ),
    .Y(_00921_));
 sky130_fd_sc_hd__inv_2 _04839_ (.A(\u_pwm.u_pwm_1.cfg_pwm_scale[0] ),
    .Y(_00922_));
 sky130_fd_sc_hd__inv_2 _04840_ (.A(\u_pwm.u_pwm_1.cfg_pwm_scale[1] ),
    .Y(_00923_));
 sky130_fd_sc_hd__inv_2 _04841_ (.A(\u_pwm.u_pwm_2.cfg_pwm_scale[2] ),
    .Y(_00924_));
 sky130_fd_sc_hd__inv_2 _04842_ (.A(\u_pwm.u_pwm_2.cfg_pwm_scale[0] ),
    .Y(_00925_));
 sky130_fd_sc_hd__inv_2 _04843_ (.A(\u_pwm.u_pwm_2.cfg_pwm_scale[1] ),
    .Y(_00926_));
 sky130_fd_sc_hd__inv_2 _04844_ (.A(\u_timer.cfg_pulse_1us[1] ),
    .Y(_00927_));
 sky130_fd_sc_hd__inv_2 _04845_ (.A(\u_timer.u_pulse_1us.cnt[3] ),
    .Y(_00928_));
 sky130_fd_sc_hd__inv_2 _04846_ (.A(\u_timer.cfg_pulse_1us[4] ),
    .Y(_00929_));
 sky130_fd_sc_hd__inv_2 _04847_ (.A(\u_timer.u_pulse_1us.cnt[6] ),
    .Y(_00930_));
 sky130_fd_sc_hd__inv_2 _04848_ (.A(\u_timer.u_pulse_1us.cnt[7] ),
    .Y(_00931_));
 sky130_fd_sc_hd__inv_2 _04849_ (.A(\u_timer.cfg_pulse_1us[7] ),
    .Y(_00932_));
 sky130_fd_sc_hd__inv_2 _04850_ (.A(\u_timer.u_pulse_1us.cnt[8] ),
    .Y(_00933_));
 sky130_fd_sc_hd__inv_2 _04851_ (.A(\u_timer.u_pulse_1us.cnt[9] ),
    .Y(_00934_));
 sky130_fd_sc_hd__inv_2 _04852_ (.A(\u_gpio.cfg_gpio_dir_sel[19] ),
    .Y(_00935_));
 sky130_fd_sc_hd__inv_2 _04853_ (.A(\u_gpio.cfg_gpio_dir_sel[18] ),
    .Y(_00936_));
 sky130_fd_sc_hd__clkinv_2 _04854_ (.A(\u_gpio.cfg_gpio_dir_sel[4] ),
    .Y(_00937_));
 sky130_fd_sc_hd__clkinv_4 _04855_ (.A(net41),
    .Y(_00938_));
 sky130_fd_sc_hd__clkinv_4 _04856_ (.A(net43),
    .Y(_00939_));
 sky130_fd_sc_hd__inv_2 _04857_ (.A(\u_gpio.cfg_gpio_dir_sel[16] ),
    .Y(net267));
 sky130_fd_sc_hd__inv_2 _04858_ (.A(\u_gpio.cfg_gpio_dir_sel[17] ),
    .Y(net268));
 sky130_fd_sc_hd__inv_2 _04859_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[14] ),
    .Y(_00940_));
 sky130_fd_sc_hd__inv_2 _04860_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[9] ),
    .Y(_00941_));
 sky130_fd_sc_hd__inv_2 _04861_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ),
    .Y(_00942_));
 sky130_fd_sc_hd__inv_2 _04862_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp0[14] ),
    .Y(_00943_));
 sky130_fd_sc_hd__inv_2 _04863_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp0[13] ),
    .Y(_00944_));
 sky130_fd_sc_hd__inv_2 _04864_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp0[10] ),
    .Y(_00945_));
 sky130_fd_sc_hd__inv_2 _04865_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[14] ),
    .Y(_00946_));
 sky130_fd_sc_hd__inv_2 _04866_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[10] ),
    .Y(_00947_));
 sky130_fd_sc_hd__inv_2 _04867_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[9] ),
    .Y(_00948_));
 sky130_fd_sc_hd__inv_2 _04868_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[8] ),
    .Y(_00949_));
 sky130_fd_sc_hd__inv_2 _04869_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[7] ),
    .Y(_00950_));
 sky130_fd_sc_hd__inv_2 _04870_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[6] ),
    .Y(_00951_));
 sky130_fd_sc_hd__inv_2 _04871_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ),
    .Y(_00952_));
 sky130_fd_sc_hd__inv_2 _04872_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ),
    .Y(_00953_));
 sky130_fd_sc_hd__inv_2 _04873_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ),
    .Y(_00954_));
 sky130_fd_sc_hd__inv_2 _04874_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ),
    .Y(_00955_));
 sky130_fd_sc_hd__inv_2 _04875_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[13] ),
    .Y(_00956_));
 sky130_fd_sc_hd__inv_2 _04876_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[10] ),
    .Y(_00957_));
 sky130_fd_sc_hd__inv_2 _04877_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[9] ),
    .Y(_00958_));
 sky130_fd_sc_hd__inv_2 _04878_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ),
    .Y(_00959_));
 sky130_fd_sc_hd__inv_2 _04879_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ),
    .Y(_00960_));
 sky130_fd_sc_hd__inv_2 _04880_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[8] ),
    .Y(_00961_));
 sky130_fd_sc_hd__inv_2 _04881_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[10] ),
    .Y(_00962_));
 sky130_fd_sc_hd__inv_2 _04882_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[11] ),
    .Y(_00963_));
 sky130_fd_sc_hd__inv_2 _04883_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ),
    .Y(_00964_));
 sky130_fd_sc_hd__inv_2 _04884_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[14] ),
    .Y(_00965_));
 sky130_fd_sc_hd__inv_2 _04885_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .Y(_00966_));
 sky130_fd_sc_hd__inv_2 _04886_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[11] ),
    .Y(_00967_));
 sky130_fd_sc_hd__inv_2 _04887_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[12] ),
    .Y(_00968_));
 sky130_fd_sc_hd__inv_2 _04888_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[13] ),
    .Y(_00969_));
 sky130_fd_sc_hd__inv_2 _04889_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[14] ),
    .Y(_00970_));
 sky130_fd_sc_hd__inv_2 _04890_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp0[14] ),
    .Y(_00971_));
 sky130_fd_sc_hd__inv_2 _04891_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ),
    .Y(_00972_));
 sky130_fd_sc_hd__inv_2 _04892_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ),
    .Y(_00973_));
 sky130_fd_sc_hd__inv_2 _04893_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ),
    .Y(_00974_));
 sky130_fd_sc_hd__inv_2 _04894_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[10] ),
    .Y(_00975_));
 sky130_fd_sc_hd__inv_2 _04895_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[9] ),
    .Y(_00976_));
 sky130_fd_sc_hd__clkinv_2 _04896_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ),
    .Y(_00977_));
 sky130_fd_sc_hd__inv_2 _04897_ (.A(\u_pwm.u_pwm_0.cfg_comp2_center ),
    .Y(_00978_));
 sky130_fd_sc_hd__inv_2 _04898_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ),
    .Y(_00979_));
 sky130_fd_sc_hd__inv_2 _04899_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[14] ),
    .Y(_00980_));
 sky130_fd_sc_hd__inv_2 _04900_ (.A(\u_pwm.u_pwm_1.cfg_comp0_center ),
    .Y(_00981_));
 sky130_fd_sc_hd__inv_2 _04901_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[0] ),
    .Y(_00982_));
 sky130_fd_sc_hd__inv_2 _04902_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[10] ),
    .Y(_00983_));
 sky130_fd_sc_hd__inv_2 _04903_ (.A(\u_pwm.u_pwm_1.cfg_comp1_center ),
    .Y(_00984_));
 sky130_fd_sc_hd__inv_2 _04904_ (.A(net1091),
    .Y(_00985_));
 sky130_fd_sc_hd__inv_2 _04905_ (.A(\reg_blk_sel[2] ),
    .Y(_00986_));
 sky130_fd_sc_hd__inv_2 _04906_ (.A(net1651),
    .Y(_00987_));
 sky130_fd_sc_hd__inv_2 _04907_ (.A(net1403),
    .Y(_00988_));
 sky130_fd_sc_hd__inv_2 _04908_ (.A(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ),
    .Y(_00989_));
 sky130_fd_sc_hd__inv_2 _04909_ (.A(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ),
    .Y(_00990_));
 sky130_fd_sc_hd__inv_2 _04910_ (.A(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ),
    .Y(_00991_));
 sky130_fd_sc_hd__or2_4 _04911_ (.A(\u_glbl_reg.cfg_gpio_dgmode ),
    .B(\u_gpio.pulse_1us ),
    .X(_00250_));
 sky130_fd_sc_hd__a31o_1 _04912_ (.A1(\u_gpio.u_bit[0].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[0].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[0].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[0].u_dglitch.gpio_reg ),
    .X(_00992_));
 sky130_fd_sc_hd__o31a_2 _04913_ (.A1(\u_gpio.u_bit[0].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[0].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[0].u_dglitch.gpio_ss[1] ),
    .B1(_00992_),
    .X(\u_gpio.u_bit[0].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _04914_ (.A_N(\u_gpio.u_bit[0].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[0] ),
    .X(_00993_));
 sky130_fd_sc_hd__and2_1 _04915_ (.A(\u_gpio.u_bit[0].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[0] ),
    .X(_00994_));
 sky130_fd_sc_hd__mux2_1 _04916_ (.A0(_00994_),
    .A1(_00993_),
    .S(\u_gpio.u_bit[0].u_dglitch.gpio_out ),
    .X(_00995_));
 sky130_fd_sc_hd__and2_2 _04917_ (.A(_00779_),
    .B(net1346),
    .X(_00996_));
 sky130_fd_sc_hd__nand2_4 _04918_ (.A(_00779_),
    .B(net1346),
    .Y(_00997_));
 sky130_fd_sc_hd__nor2_1 _04919_ (.A(net1358),
    .B(net1264),
    .Y(_00998_));
 sky130_fd_sc_hd__nand2_8 _04920_ (.A(net1267),
    .B(net1362),
    .Y(_00999_));
 sky130_fd_sc_hd__nor2_4 _04921_ (.A(net1359),
    .B(_00997_),
    .Y(_01000_));
 sky130_fd_sc_hd__nor2_2 _04922_ (.A(_00997_),
    .B(_00999_),
    .Y(_01001_));
 sky130_fd_sc_hd__and2b_2 _04923_ (.A_N(net1341),
    .B(net1307),
    .X(_01002_));
 sky130_fd_sc_hd__nor2_2 _04924_ (.A(net1374),
    .B(net1340),
    .Y(_01003_));
 sky130_fd_sc_hd__and4_1 _04925_ (.A(net1416),
    .B(net1342),
    .C(_01002_),
    .D(_01003_),
    .X(_01004_));
 sky130_fd_sc_hd__and3_2 _04926_ (.A(\u_gpio.reg_ack ),
    .B(_01001_),
    .C(net1177),
    .X(_01005_));
 sky130_fd_sc_hd__a21o_1 _04927_ (.A1(net1296),
    .A2(net577),
    .B1(_00995_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__nor2_1 _04928_ (.A(net1359),
    .B(net1368),
    .Y(_01006_));
 sky130_fd_sc_hd__or2_1 _04929_ (.A(net1356),
    .B(net1364),
    .X(_01007_));
 sky130_fd_sc_hd__nor2_1 _04930_ (.A(_00997_),
    .B(net1228),
    .Y(_01008_));
 sky130_fd_sc_hd__a41o_4 _04931_ (.A1(\u_gpio.reg_ack ),
    .A2(net1336),
    .A3(net1177),
    .A4(net711),
    .B1(net577),
    .X(_01009_));
 sky130_fd_sc_hd__a21o_1 _04932_ (.A1(net1296),
    .A2(_01009_),
    .B1(_00995_),
    .X(_00264_));
 sky130_fd_sc_hd__a31o_1 _04933_ (.A1(\u_gpio.u_bit[10].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[10].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[10].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[10].u_dglitch.gpio_reg ),
    .X(_01010_));
 sky130_fd_sc_hd__o31a_1 _04934_ (.A1(\u_gpio.u_bit[10].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[10].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[10].u_dglitch.gpio_ss[1] ),
    .B1(_01010_),
    .X(\u_gpio.u_bit[10].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04935_ (.A(\u_gpio.u_bit[10].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[10] ),
    .Y(_01011_));
 sky130_fd_sc_hd__a2bb2o_1 _04936_ (.A1_N(\u_gpio.u_bit[10].u_dglitch.gpio_out ),
    .A2_N(_01011_),
    .B1(net1286),
    .B2(net576),
    .X(_01012_));
 sky130_fd_sc_hd__a31o_1 _04937_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[10] ),
    .A2(_00780_),
    .A3(\u_gpio.u_bit[10].u_dglitch.gpio_out ),
    .B1(_01012_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and4_4 _04938_ (.A(\u_gpio.reg_ack ),
    .B(net1327),
    .C(net1177),
    .D(net711),
    .X(_01013_));
 sky130_fd_sc_hd__a21o_1 _04939_ (.A1(net1287),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.hware_req ),
    .X(_00265_));
 sky130_fd_sc_hd__a31o_1 _04940_ (.A1(\u_gpio.u_bit[11].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[11].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[11].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[11].u_dglitch.gpio_reg ),
    .X(_01014_));
 sky130_fd_sc_hd__o31a_1 _04941_ (.A1(\u_gpio.u_bit[11].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[11].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[11].u_dglitch.gpio_ss[1] ),
    .B1(_01014_),
    .X(\u_gpio.u_bit[11].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04942_ (.A(\u_gpio.u_bit[11].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[11] ),
    .Y(_01015_));
 sky130_fd_sc_hd__a2bb2o_1 _04943_ (.A1_N(\u_gpio.u_bit[11].u_dglitch.gpio_out ),
    .A2_N(_01015_),
    .B1(net1643),
    .B2(net576),
    .X(_01016_));
 sky130_fd_sc_hd__a31o_1 _04944_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[11] ),
    .A2(_00781_),
    .A3(\u_gpio.u_bit[11].u_dglitch.gpio_out ),
    .B1(_01016_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04945_ (.A1(net1643),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.hware_req ),
    .X(_00266_));
 sky130_fd_sc_hd__a31o_1 _04946_ (.A1(\u_gpio.u_bit[12].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[12].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[12].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[12].u_dglitch.gpio_reg ),
    .X(_01017_));
 sky130_fd_sc_hd__o31a_1 _04947_ (.A1(\u_gpio.u_bit[12].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[12].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[12].u_dglitch.gpio_ss[1] ),
    .B1(_01017_),
    .X(\u_gpio.u_bit[12].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04948_ (.A(\u_gpio.u_bit[12].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[12] ),
    .Y(_01018_));
 sky130_fd_sc_hd__a2bb2o_1 _04949_ (.A1_N(\u_gpio.u_bit[12].u_dglitch.gpio_out ),
    .A2_N(_01018_),
    .B1(net1636),
    .B2(net575),
    .X(_01019_));
 sky130_fd_sc_hd__a31o_1 _04950_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[12] ),
    .A2(_00782_),
    .A3(\u_gpio.u_bit[12].u_dglitch.gpio_out ),
    .B1(_01019_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04951_ (.A1(net1636),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.hware_req ),
    .X(_00267_));
 sky130_fd_sc_hd__a31o_1 _04952_ (.A1(\u_gpio.u_bit[13].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[13].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[13].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[13].u_dglitch.gpio_reg ),
    .X(_01020_));
 sky130_fd_sc_hd__o31a_1 _04953_ (.A1(\u_gpio.u_bit[13].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[13].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[13].u_dglitch.gpio_ss[1] ),
    .B1(_01020_),
    .X(\u_gpio.u_bit[13].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04954_ (.A(\u_gpio.u_bit[13].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[13] ),
    .Y(_01021_));
 sky130_fd_sc_hd__a2bb2o_1 _04955_ (.A1_N(\u_gpio.u_bit[13].u_dglitch.gpio_out ),
    .A2_N(_01021_),
    .B1(net1628),
    .B2(net577),
    .X(_01022_));
 sky130_fd_sc_hd__a31o_1 _04956_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[13] ),
    .A2(_00783_),
    .A3(\u_gpio.u_bit[13].u_dglitch.gpio_out ),
    .B1(_01022_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04957_ (.A1(net1628),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.hware_req ),
    .X(_00268_));
 sky130_fd_sc_hd__a31o_1 _04958_ (.A1(\u_gpio.u_bit[14].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[14].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[14].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[14].u_dglitch.gpio_reg ),
    .X(_01023_));
 sky130_fd_sc_hd__o31a_1 _04959_ (.A1(\u_gpio.u_bit[14].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[14].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[14].u_dglitch.gpio_ss[1] ),
    .B1(_01023_),
    .X(\u_gpio.u_bit[14].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04960_ (.A(\u_gpio.u_bit[14].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[14] ),
    .Y(_01024_));
 sky130_fd_sc_hd__a2bb2o_1 _04961_ (.A1_N(\u_gpio.u_bit[14].u_dglitch.gpio_out ),
    .A2_N(_01024_),
    .B1(net1621),
    .B2(net577),
    .X(_01025_));
 sky130_fd_sc_hd__a31o_1 _04962_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[14] ),
    .A2(_00784_),
    .A3(\u_gpio.u_bit[14].u_dglitch.gpio_out ),
    .B1(_01025_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04963_ (.A1(net1621),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.hware_req ),
    .X(_00269_));
 sky130_fd_sc_hd__a31o_1 _04964_ (.A1(\u_gpio.u_bit[15].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[15].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[15].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[15].u_dglitch.gpio_reg ),
    .X(_01026_));
 sky130_fd_sc_hd__o31a_1 _04965_ (.A1(\u_gpio.u_bit[15].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[15].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[15].u_dglitch.gpio_ss[1] ),
    .B1(_01026_),
    .X(\u_gpio.u_bit[15].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _04966_ (.A(\u_gpio.u_bit[15].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[15] ),
    .Y(_01027_));
 sky130_fd_sc_hd__a2bb2o_1 _04967_ (.A1_N(\u_gpio.u_bit[15].u_dglitch.gpio_out ),
    .A2_N(_01027_),
    .B1(net1615),
    .B2(net577),
    .X(_01028_));
 sky130_fd_sc_hd__a31o_1 _04968_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[15] ),
    .A2(_00785_),
    .A3(\u_gpio.u_bit[15].u_dglitch.gpio_out ),
    .B1(_01028_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04969_ (.A1(net1615),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.hware_req ),
    .X(_00270_));
 sky130_fd_sc_hd__a31o_1 _04970_ (.A1(\u_gpio.u_bit[16].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[16].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[16].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[16].u_dglitch.gpio_reg ),
    .X(_01029_));
 sky130_fd_sc_hd__o31a_4 _04971_ (.A1(\u_gpio.u_bit[16].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[16].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[16].u_dglitch.gpio_ss[1] ),
    .B1(_01029_),
    .X(\u_gpio.u_bit[16].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _04972_ (.A_N(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[16] ),
    .C(\u_gpio.u_bit[16].u_dglitch.gpio_reg ),
    .X(_01030_));
 sky130_fd_sc_hd__a31o_1 _04973_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[16] ),
    .A2(_00786_),
    .A3(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .B1(_01030_),
    .X(_01031_));
 sky130_fd_sc_hd__a21o_1 _04974_ (.A1(net1607),
    .A2(net578),
    .B1(_01031_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a41o_1 _04975_ (.A1(\u_gpio.reg_ack ),
    .A2(net1318),
    .A3(net1177),
    .A4(net711),
    .B1(net577),
    .X(_01032_));
 sky130_fd_sc_hd__a21o_1 _04976_ (.A1(net1607),
    .A2(net535),
    .B1(_01031_),
    .X(_00271_));
 sky130_fd_sc_hd__a31o_1 _04977_ (.A1(\u_gpio.u_bit[17].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[17].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[17].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[17].u_dglitch.gpio_reg ),
    .X(_01033_));
 sky130_fd_sc_hd__o31a_4 _04978_ (.A1(\u_gpio.u_bit[17].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[17].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[17].u_dglitch.gpio_ss[1] ),
    .B1(_01033_),
    .X(\u_gpio.u_bit[17].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _04979_ (.A_N(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[17] ),
    .C(\u_gpio.u_bit[17].u_dglitch.gpio_reg ),
    .X(_01034_));
 sky130_fd_sc_hd__a31o_1 _04980_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[17] ),
    .A2(_00787_),
    .A3(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .B1(_01034_),
    .X(_01035_));
 sky130_fd_sc_hd__a21o_1 _04981_ (.A1(net1600),
    .A2(net578),
    .B1(_01035_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04982_ (.A1(net1600),
    .A2(net535),
    .B1(_01035_),
    .X(_00272_));
 sky130_fd_sc_hd__a31o_1 _04983_ (.A1(\u_gpio.u_bit[18].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[18].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[18].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[18].u_dglitch.gpio_reg ),
    .X(_01036_));
 sky130_fd_sc_hd__o31a_4 _04984_ (.A1(\u_gpio.u_bit[18].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[18].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[18].u_dglitch.gpio_ss[1] ),
    .B1(_01036_),
    .X(\u_gpio.u_bit[18].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _04985_ (.A_N(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[18] ),
    .C(\u_gpio.u_bit[18].u_dglitch.gpio_reg ),
    .X(_01037_));
 sky130_fd_sc_hd__a31o_1 _04986_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[18] ),
    .A2(_00788_),
    .A3(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .B1(_01037_),
    .X(_01038_));
 sky130_fd_sc_hd__a21o_1 _04987_ (.A1(net1586),
    .A2(net578),
    .B1(_01038_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04988_ (.A1(net1587),
    .A2(net535),
    .B1(_01038_),
    .X(_00273_));
 sky130_fd_sc_hd__a31o_1 _04989_ (.A1(\u_gpio.u_bit[19].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[19].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[19].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[19].u_dglitch.gpio_reg ),
    .X(_01039_));
 sky130_fd_sc_hd__o31ai_4 _04990_ (.A1(\u_gpio.u_bit[19].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[19].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[19].u_dglitch.gpio_ss[1] ),
    .B1(_01039_),
    .Y(_01040_));
 sky130_fd_sc_hd__inv_2 _04991_ (.A(_01040_),
    .Y(\u_gpio.u_bit[19].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _04992_ (.A_N(\u_gpio.u_bit[19].u_dglitch.gpio_reg ),
    .B(\u_gpio.u_bit[19].u_dglitch.gpio_out ),
    .C(\u_gpio.cfg_gpio_posedge_int_sel[19] ),
    .X(_01041_));
 sky130_fd_sc_hd__a31o_1 _04993_ (.A1(\u_gpio.u_bit[19].u_dglitch.gpio_reg ),
    .A2(\u_gpio.cfg_gpio_negedge_int_sel[19] ),
    .A3(_01040_),
    .B1(_01041_),
    .X(_01042_));
 sky130_fd_sc_hd__a21o_1 _04994_ (.A1(net1581),
    .A2(net578),
    .B1(_01042_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _04995_ (.A1(net1581),
    .A2(net535),
    .B1(_01042_),
    .X(_00274_));
 sky130_fd_sc_hd__a31o_1 _04996_ (.A1(\u_gpio.u_bit[1].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[1].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[1].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[1].u_dglitch.gpio_reg ),
    .X(_01043_));
 sky130_fd_sc_hd__o31a_1 _04997_ (.A1(\u_gpio.u_bit[1].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[1].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[1].u_dglitch.gpio_ss[1] ),
    .B1(_01043_),
    .X(\u_gpio.u_bit[1].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _04998_ (.A_N(\u_gpio.u_bit[1].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[1] ),
    .X(_01044_));
 sky130_fd_sc_hd__and2_1 _04999_ (.A(\u_gpio.u_bit[1].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[1] ),
    .X(_01045_));
 sky130_fd_sc_hd__mux2_1 _05000_ (.A0(_01045_),
    .A1(_01044_),
    .S(\u_gpio.u_bit[1].u_dglitch.gpio_out ),
    .X(_01046_));
 sky130_fd_sc_hd__a21o_1 _05001_ (.A1(net1575),
    .A2(net576),
    .B1(_01046_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05002_ (.A1(net1575),
    .A2(_01009_),
    .B1(_01046_),
    .X(_00275_));
 sky130_fd_sc_hd__a31o_1 _05003_ (.A1(\u_gpio.u_bit[20].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[20].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[20].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[20].u_dglitch.gpio_reg ),
    .X(_01047_));
 sky130_fd_sc_hd__o31a_4 _05004_ (.A1(\u_gpio.u_bit[20].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[20].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[20].u_dglitch.gpio_ss[1] ),
    .B1(_01047_),
    .X(\u_gpio.u_bit[20].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _05005_ (.A_N(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[20] ),
    .C(\u_gpio.u_bit[20].u_dglitch.gpio_reg ),
    .X(_01048_));
 sky130_fd_sc_hd__a31o_1 _05006_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[20] ),
    .A2(_00789_),
    .A3(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .B1(_01048_),
    .X(_01049_));
 sky130_fd_sc_hd__a21o_1 _05007_ (.A1(net1566),
    .A2(net578),
    .B1(_01049_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05008_ (.A1(net1566),
    .A2(net535),
    .B1(_01049_),
    .X(_00276_));
 sky130_fd_sc_hd__a31o_1 _05009_ (.A1(\u_gpio.u_bit[21].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[21].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[21].u_dglitch.gpio_reg ),
    .X(_01050_));
 sky130_fd_sc_hd__o31a_4 _05010_ (.A1(\u_gpio.u_bit[21].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[21].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_ss[1] ),
    .B1(_01050_),
    .X(\u_gpio.u_bit[21].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _05011_ (.A_N(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[21] ),
    .C(\u_gpio.u_bit[21].u_dglitch.gpio_reg ),
    .X(_01051_));
 sky130_fd_sc_hd__a31o_1 _05012_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[21] ),
    .A2(_00790_),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .B1(_01051_),
    .X(_01052_));
 sky130_fd_sc_hd__a21o_1 _05013_ (.A1(net1559),
    .A2(net578),
    .B1(_01052_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05014_ (.A1(net1559),
    .A2(net535),
    .B1(_01052_),
    .X(_00277_));
 sky130_fd_sc_hd__a31o_1 _05015_ (.A1(\u_gpio.u_bit[22].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[22].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[22].u_dglitch.gpio_reg ),
    .X(_01053_));
 sky130_fd_sc_hd__o31a_4 _05016_ (.A1(\u_gpio.u_bit[22].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[22].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_ss[1] ),
    .B1(_01053_),
    .X(\u_gpio.u_bit[22].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and3b_1 _05017_ (.A_N(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[22] ),
    .C(\u_gpio.u_bit[22].u_dglitch.gpio_reg ),
    .X(_01054_));
 sky130_fd_sc_hd__a31o_1 _05018_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[22] ),
    .A2(_00791_),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .B1(_01054_),
    .X(_01055_));
 sky130_fd_sc_hd__a21o_1 _05019_ (.A1(net1551),
    .A2(net577),
    .B1(_01055_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05020_ (.A1(net1551),
    .A2(net534),
    .B1(_01055_),
    .X(_00278_));
 sky130_fd_sc_hd__and2_1 _05021_ (.A(net1542),
    .B(net578),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_1 _05022_ (.A(net1542),
    .B(net534),
    .X(_00279_));
 sky130_fd_sc_hd__a31o_1 _05023_ (.A1(\u_gpio.u_bit[24].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[24].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[24].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[24].u_dglitch.gpio_reg ),
    .X(_01056_));
 sky130_fd_sc_hd__o31a_1 _05024_ (.A1(\u_gpio.u_bit[24].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[24].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[24].u_dglitch.gpio_ss[1] ),
    .B1(_01056_),
    .X(\u_gpio.u_bit[24].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05025_ (.A_N(\u_gpio.u_bit[24].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[24] ),
    .X(_01057_));
 sky130_fd_sc_hd__and2_1 _05026_ (.A(\u_gpio.u_bit[24].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[24] ),
    .X(_01058_));
 sky130_fd_sc_hd__mux2_1 _05027_ (.A0(_01058_),
    .A1(_01057_),
    .S(\u_gpio.u_bit[24].u_dglitch.gpio_out ),
    .X(_01059_));
 sky130_fd_sc_hd__a21o_1 _05028_ (.A1(net1536),
    .A2(net575),
    .B1(_01059_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05029_ (.A1(net1536),
    .A2(net534),
    .B1(_01059_),
    .X(_00280_));
 sky130_fd_sc_hd__a31o_1 _05030_ (.A1(\u_gpio.u_bit[25].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[25].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[25].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[25].u_dglitch.gpio_reg ),
    .X(_01060_));
 sky130_fd_sc_hd__o31a_2 _05031_ (.A1(\u_gpio.u_bit[25].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[25].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[25].u_dglitch.gpio_ss[1] ),
    .B1(_01060_),
    .X(\u_gpio.u_bit[25].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05032_ (.A_N(\u_gpio.u_bit[25].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[25] ),
    .X(_01061_));
 sky130_fd_sc_hd__and2_1 _05033_ (.A(\u_gpio.u_bit[25].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[25] ),
    .X(_01062_));
 sky130_fd_sc_hd__mux2_1 _05034_ (.A0(_01062_),
    .A1(_01061_),
    .S(\u_gpio.u_bit[25].u_dglitch.gpio_out ),
    .X(_01063_));
 sky130_fd_sc_hd__a21o_1 _05035_ (.A1(net1528),
    .A2(net575),
    .B1(_01063_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05036_ (.A1(net1528),
    .A2(net534),
    .B1(_01063_),
    .X(_00281_));
 sky130_fd_sc_hd__a31o_1 _05037_ (.A1(\u_gpio.u_bit[26].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[26].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[26].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[26].u_dglitch.gpio_reg ),
    .X(_01064_));
 sky130_fd_sc_hd__o31a_1 _05038_ (.A1(\u_gpio.u_bit[26].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[26].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[26].u_dglitch.gpio_ss[1] ),
    .B1(_01064_),
    .X(\u_gpio.u_bit[26].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05039_ (.A_N(\u_gpio.u_bit[26].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[26] ),
    .X(_01065_));
 sky130_fd_sc_hd__and2_1 _05040_ (.A(\u_gpio.u_bit[26].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[26] ),
    .X(_01066_));
 sky130_fd_sc_hd__mux2_1 _05041_ (.A0(_01066_),
    .A1(_01065_),
    .S(\u_gpio.u_bit[26].u_dglitch.gpio_out ),
    .X(_01067_));
 sky130_fd_sc_hd__a21o_1 _05042_ (.A1(net1521),
    .A2(net575),
    .B1(_01067_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05043_ (.A1(net1521),
    .A2(net534),
    .B1(_01067_),
    .X(_00282_));
 sky130_fd_sc_hd__a31o_1 _05044_ (.A1(\u_gpio.u_bit[27].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[27].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[27].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[27].u_dglitch.gpio_reg ),
    .X(_01068_));
 sky130_fd_sc_hd__o31a_2 _05045_ (.A1(\u_gpio.u_bit[27].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[27].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[27].u_dglitch.gpio_ss[1] ),
    .B1(_01068_),
    .X(\u_gpio.u_bit[27].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05046_ (.A_N(\u_gpio.u_bit[27].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[27] ),
    .X(_01069_));
 sky130_fd_sc_hd__and2_1 _05047_ (.A(\u_gpio.u_bit[27].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[27] ),
    .X(_01070_));
 sky130_fd_sc_hd__mux2_1 _05048_ (.A0(_01070_),
    .A1(_01069_),
    .S(\u_gpio.u_bit[27].u_dglitch.gpio_out ),
    .X(_01071_));
 sky130_fd_sc_hd__a21o_1 _05049_ (.A1(net1514),
    .A2(net575),
    .B1(_01071_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05050_ (.A1(net1514),
    .A2(net534),
    .B1(_01071_),
    .X(_00283_));
 sky130_fd_sc_hd__a31o_1 _05051_ (.A1(\u_gpio.u_bit[28].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[28].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[28].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[28].u_dglitch.gpio_reg ),
    .X(_01072_));
 sky130_fd_sc_hd__o31a_2 _05052_ (.A1(\u_gpio.u_bit[28].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[28].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[28].u_dglitch.gpio_ss[1] ),
    .B1(_01072_),
    .X(\u_gpio.u_bit[28].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05053_ (.A_N(\u_gpio.u_bit[28].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[28] ),
    .X(_01073_));
 sky130_fd_sc_hd__and2_1 _05054_ (.A(\u_gpio.u_bit[28].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[28] ),
    .X(_01074_));
 sky130_fd_sc_hd__mux2_1 _05055_ (.A0(_01074_),
    .A1(_01073_),
    .S(\u_gpio.u_bit[28].u_dglitch.gpio_out ),
    .X(_01075_));
 sky130_fd_sc_hd__a21o_1 _05056_ (.A1(net1508),
    .A2(net575),
    .B1(_01075_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05057_ (.A1(net1508),
    .A2(net534),
    .B1(_01075_),
    .X(_00284_));
 sky130_fd_sc_hd__a31o_1 _05058_ (.A1(\u_gpio.u_bit[29].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[29].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[29].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[29].u_dglitch.gpio_reg ),
    .X(_01076_));
 sky130_fd_sc_hd__o31a_1 _05059_ (.A1(\u_gpio.u_bit[29].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[29].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[29].u_dglitch.gpio_ss[1] ),
    .B1(_01076_),
    .X(\u_gpio.u_bit[29].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05060_ (.A_N(\u_gpio.u_bit[29].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[29] ),
    .X(_01077_));
 sky130_fd_sc_hd__and2_1 _05061_ (.A(\u_gpio.u_bit[29].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[29] ),
    .X(_01078_));
 sky130_fd_sc_hd__mux2_1 _05062_ (.A0(_01078_),
    .A1(_01077_),
    .S(\u_gpio.u_bit[29].u_dglitch.gpio_out ),
    .X(_01079_));
 sky130_fd_sc_hd__a21o_1 _05063_ (.A1(net1499),
    .A2(net575),
    .B1(_01079_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05064_ (.A1(net1499),
    .A2(net534),
    .B1(_01079_),
    .X(_00285_));
 sky130_fd_sc_hd__a31o_1 _05065_ (.A1(\u_gpio.u_bit[2].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[2].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[2].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[2].u_dglitch.gpio_reg ),
    .X(_01080_));
 sky130_fd_sc_hd__o31a_1 _05066_ (.A1(\u_gpio.u_bit[2].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[2].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[2].u_dglitch.gpio_ss[1] ),
    .B1(_01080_),
    .X(\u_gpio.u_bit[2].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05067_ (.A_N(\u_gpio.u_bit[2].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[2] ),
    .X(_01081_));
 sky130_fd_sc_hd__and2_1 _05068_ (.A(\u_gpio.u_bit[2].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[2] ),
    .X(_01082_));
 sky130_fd_sc_hd__mux2_1 _05069_ (.A0(_01082_),
    .A1(_01081_),
    .S(\u_gpio.u_bit[2].u_dglitch.gpio_out ),
    .X(_01083_));
 sky130_fd_sc_hd__a21o_1 _05070_ (.A1(net1490),
    .A2(net577),
    .B1(_01083_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05071_ (.A1(net1490),
    .A2(_01009_),
    .B1(_01083_),
    .X(_00286_));
 sky130_fd_sc_hd__a31o_1 _05072_ (.A1(\u_gpio.u_bit[30].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[30].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[30].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[30].u_dglitch.gpio_reg ),
    .X(_01084_));
 sky130_fd_sc_hd__o31a_1 _05073_ (.A1(\u_gpio.u_bit[30].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[30].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[30].u_dglitch.gpio_ss[1] ),
    .B1(_01084_),
    .X(\u_gpio.u_bit[30].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05074_ (.A_N(\u_gpio.u_bit[30].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[30] ),
    .X(_01085_));
 sky130_fd_sc_hd__and2_1 _05075_ (.A(\u_gpio.u_bit[30].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[30] ),
    .X(_01086_));
 sky130_fd_sc_hd__mux2_1 _05076_ (.A0(_01086_),
    .A1(_01085_),
    .S(\u_gpio.u_bit[30].u_dglitch.gpio_out ),
    .X(_01087_));
 sky130_fd_sc_hd__a21o_1 _05077_ (.A1(net1483),
    .A2(net575),
    .B1(_01087_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05078_ (.A1(net1483),
    .A2(net534),
    .B1(_01087_),
    .X(_00287_));
 sky130_fd_sc_hd__a31o_1 _05079_ (.A1(\u_gpio.u_bit[31].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[31].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[31].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[31].u_dglitch.gpio_reg ),
    .X(_01088_));
 sky130_fd_sc_hd__o31a_1 _05080_ (.A1(\u_gpio.u_bit[31].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[31].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[31].u_dglitch.gpio_ss[1] ),
    .B1(_01088_),
    .X(\u_gpio.u_bit[31].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05081_ (.A_N(\u_gpio.u_bit[31].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[31] ),
    .X(_01089_));
 sky130_fd_sc_hd__and2_1 _05082_ (.A(\u_gpio.u_bit[31].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[31] ),
    .X(_01090_));
 sky130_fd_sc_hd__mux2_1 _05083_ (.A0(_01090_),
    .A1(_01089_),
    .S(\u_gpio.u_bit[31].u_dglitch.gpio_out ),
    .X(_01091_));
 sky130_fd_sc_hd__a21o_1 _05084_ (.A1(net1476),
    .A2(net575),
    .B1(_01091_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05085_ (.A1(net1476),
    .A2(net534),
    .B1(_01091_),
    .X(_00288_));
 sky130_fd_sc_hd__a31o_1 _05086_ (.A1(\u_gpio.u_bit[3].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[3].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[3].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[3].u_dglitch.gpio_reg ),
    .X(_01092_));
 sky130_fd_sc_hd__o31a_1 _05087_ (.A1(\u_gpio.u_bit[3].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[3].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[3].u_dglitch.gpio_ss[1] ),
    .B1(_01092_),
    .X(\u_gpio.u_bit[3].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05088_ (.A_N(\u_gpio.u_bit[3].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[3] ),
    .X(_01093_));
 sky130_fd_sc_hd__and2_1 _05089_ (.A(\u_gpio.u_bit[3].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[3] ),
    .X(_01094_));
 sky130_fd_sc_hd__mux2_1 _05090_ (.A0(_01094_),
    .A1(_01093_),
    .S(\u_gpio.u_bit[3].u_dglitch.gpio_out ),
    .X(_01095_));
 sky130_fd_sc_hd__a21o_1 _05091_ (.A1(net1467),
    .A2(net576),
    .B1(_01095_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05092_ (.A1(net1467),
    .A2(_01009_),
    .B1(_01095_),
    .X(_00289_));
 sky130_fd_sc_hd__a31o_1 _05093_ (.A1(\u_gpio.u_bit[4].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[4].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[4].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[4].u_dglitch.gpio_reg ),
    .X(_01096_));
 sky130_fd_sc_hd__o31a_2 _05094_ (.A1(\u_gpio.u_bit[4].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[4].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[4].u_dglitch.gpio_ss[1] ),
    .B1(_01096_),
    .X(\u_gpio.u_bit[4].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__and2b_1 _05095_ (.A_N(\u_gpio.u_bit[4].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_posedge_int_sel[4] ),
    .X(_01097_));
 sky130_fd_sc_hd__and2_1 _05096_ (.A(\u_gpio.u_bit[4].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[4] ),
    .X(_01098_));
 sky130_fd_sc_hd__mux2_1 _05097_ (.A0(_01098_),
    .A1(_01097_),
    .S(\u_gpio.u_bit[4].u_dglitch.gpio_out ),
    .X(_01099_));
 sky130_fd_sc_hd__a21o_1 _05098_ (.A1(net1460),
    .A2(net576),
    .B1(_01099_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05099_ (.A1(net1460),
    .A2(_01009_),
    .B1(_01099_),
    .X(_00290_));
 sky130_fd_sc_hd__and2_1 _05100_ (.A(net1450),
    .B(net577),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_1 _05101_ (.A(net1450),
    .B(_01009_),
    .X(_00291_));
 sky130_fd_sc_hd__and2_1 _05102_ (.A(net1444),
    .B(net578),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_1 _05103_ (.A(net1444),
    .B(_01009_),
    .X(_00292_));
 sky130_fd_sc_hd__and2_1 _05104_ (.A(net1436),
    .B(net576),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_1 _05105_ (.A(net1436),
    .B(_01009_),
    .X(_00293_));
 sky130_fd_sc_hd__a31o_1 _05106_ (.A1(\u_gpio.u_bit[8].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[8].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[8].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[8].u_dglitch.gpio_reg ),
    .X(_01100_));
 sky130_fd_sc_hd__o31a_1 _05107_ (.A1(\u_gpio.u_bit[8].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[8].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[8].u_dglitch.gpio_ss[1] ),
    .B1(_01100_),
    .X(\u_gpio.u_bit[8].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _05108_ (.A(\u_gpio.u_bit[8].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[8] ),
    .Y(_01101_));
 sky130_fd_sc_hd__a2bb2o_1 _05109_ (.A1_N(\u_gpio.u_bit[8].u_dglitch.gpio_out ),
    .A2_N(_01101_),
    .B1(net1426),
    .B2(net577),
    .X(_01102_));
 sky130_fd_sc_hd__a31o_1 _05110_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[8] ),
    .A2(_00792_),
    .A3(\u_gpio.u_bit[8].u_dglitch.gpio_out ),
    .B1(_01102_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05111_ (.A1(net1426),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.hware_req ),
    .X(_00294_));
 sky130_fd_sc_hd__a31o_1 _05112_ (.A1(\u_gpio.u_bit[9].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[9].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[9].u_dglitch.gpio_ss[1] ),
    .B1(\u_gpio.u_bit[9].u_dglitch.gpio_reg ),
    .X(_01103_));
 sky130_fd_sc_hd__o31a_1 _05113_ (.A1(\u_gpio.u_bit[9].u_dglitch.gpio_ss[2] ),
    .A2(\u_gpio.u_bit[9].u_dglitch.gpio_ss[3] ),
    .A3(\u_gpio.u_bit[9].u_dglitch.gpio_ss[1] ),
    .B1(_01103_),
    .X(\u_gpio.u_bit[9].u_dglitch.gpio_out ));
 sky130_fd_sc_hd__nand2_1 _05114_ (.A(\u_gpio.u_bit[9].u_dglitch.gpio_reg ),
    .B(\u_gpio.cfg_gpio_negedge_int_sel[9] ),
    .Y(_01104_));
 sky130_fd_sc_hd__a2bb2o_1 _05115_ (.A1_N(\u_gpio.u_bit[9].u_dglitch.gpio_out ),
    .A2_N(_01104_),
    .B1(net1420),
    .B2(net575),
    .X(_01105_));
 sky130_fd_sc_hd__a31o_1 _05116_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[9] ),
    .A2(_00793_),
    .A3(\u_gpio.u_bit[9].u_dglitch.gpio_out ),
    .B1(_01105_),
    .X(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05117_ (.A1(net1420),
    .A2(_01013_),
    .B1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.hware_req ),
    .X(_00295_));
 sky130_fd_sc_hd__or3_1 _05118_ (.A(\u_glbl_reg.u_dbgclk.high_count[1] ),
    .B(\u_glbl_reg.u_dbgclk.high_count[0] ),
    .C(\u_glbl_reg.u_dbgclk.high_count[2] ),
    .X(_01106_));
 sky130_fd_sc_hd__nor2_1 _05119_ (.A(\u_glbl_reg.u_dbgclk.high_count[3] ),
    .B(_01106_),
    .Y(_00045_));
 sky130_fd_sc_hd__or2_1 _05120_ (.A(\u_glbl_reg.u_dbgclk.low_count[0] ),
    .B(\u_glbl_reg.u_dbgclk.low_count[1] ),
    .X(_01107_));
 sky130_fd_sc_hd__or3_1 _05121_ (.A(\u_glbl_reg.u_dbgclk.low_count[3] ),
    .B(\u_glbl_reg.u_dbgclk.low_count[2] ),
    .C(_01107_),
    .X(_01108_));
 sky130_fd_sc_hd__nand2_1 _05122_ (.A(_00045_),
    .B(_01108_),
    .Y(_00044_));
 sky130_fd_sc_hd__or2_1 _05123_ (.A(\u_glbl_reg.u_pll_ref_clk.high_count[1] ),
    .B(\u_glbl_reg.u_pll_ref_clk.high_count[0] ),
    .X(_01109_));
 sky130_fd_sc_hd__nor2_1 _05124_ (.A(\u_glbl_reg.u_pll_ref_clk.high_count[2] ),
    .B(_01109_),
    .Y(_00055_));
 sky130_fd_sc_hd__or2_1 _05125_ (.A(\u_glbl_reg.u_pll_ref_clk.low_count[0] ),
    .B(\u_glbl_reg.u_pll_ref_clk.low_count[1] ),
    .X(_01110_));
 sky130_fd_sc_hd__nor2_1 _05126_ (.A(\u_glbl_reg.u_pll_ref_clk.low_count[2] ),
    .B(_01110_),
    .Y(_01111_));
 sky130_fd_sc_hd__or2_1 _05127_ (.A(\u_glbl_reg.u_pll_ref_clk.low_count[2] ),
    .B(_01110_),
    .X(_01112_));
 sky130_fd_sc_hd__nand2_1 _05128_ (.A(_00055_),
    .B(_01112_),
    .Y(_00054_));
 sky130_fd_sc_hd__and4b_2 _05129_ (.A_N(net1342),
    .B(_01002_),
    .C(_01003_),
    .D(net1416),
    .X(_01113_));
 sky130_fd_sc_hd__nor2_8 _05130_ (.A(net1271),
    .B(net1364),
    .Y(_01114_));
 sky130_fd_sc_hd__nand2_8 _05131_ (.A(net1356),
    .B(net1260),
    .Y(_01115_));
 sky130_fd_sc_hd__nor2_1 _05132_ (.A(_00779_),
    .B(net1346),
    .Y(_01116_));
 sky130_fd_sc_hd__or2_1 _05133_ (.A(_00779_),
    .B(net1346),
    .X(_01117_));
 sky130_fd_sc_hd__nor2_4 _05134_ (.A(net1344),
    .B(_01117_),
    .Y(_01118_));
 sky130_fd_sc_hd__and4_4 _05135_ (.A(\u_glbl_reg.reg_ack ),
    .B(net1172),
    .C(net1161),
    .D(_01118_),
    .X(_01119_));
 sky130_fd_sc_hd__and2_2 _05136_ (.A(net1323),
    .B(_01119_),
    .X(_01120_));
 sky130_fd_sc_hd__a22o_1 _05137_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[9] ),
    .A2(net2304),
    .B1(_01120_),
    .B2(net1420),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and4_2 _05138_ (.A(\u_glbl_reg.reg_ack ),
    .B(net1254),
    .C(net711),
    .D(net1172),
    .X(_01121_));
 sky130_fd_sc_hd__and2_2 _05139_ (.A(net1325),
    .B(_01121_),
    .X(_01122_));
 sky130_fd_sc_hd__a21o_1 _05140_ (.A1(net1420),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.hware_req ),
    .X(_00090_));
 sky130_fd_sc_hd__a22o_1 _05141_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[8] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1426),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05142_ (.A1(net1425),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.hware_req ),
    .X(_00089_));
 sky130_fd_sc_hd__and2_4 _05143_ (.A(net1336),
    .B(_01119_),
    .X(_01123_));
 sky130_fd_sc_hd__a31o_1 _05144_ (.A1(net1336),
    .A2(net1438),
    .A3(_01119_),
    .B1(\u_glbl_reg.ir_intr_ss ),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_4 _05145_ (.A(net1335),
    .B(_01121_),
    .X(_01124_));
 sky130_fd_sc_hd__a21o_1 _05146_ (.A1(net1438),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.hware_req ),
    .X(_00088_));
 sky130_fd_sc_hd__a31o_1 _05147_ (.A1(net1336),
    .A2(net1447),
    .A3(_01119_),
    .B1(\u_glbl_reg.rtc_intr_ss ),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05148_ (.A1(net1445),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.hware_req ),
    .X(_00087_));
 sky130_fd_sc_hd__and2_2 _05149_ (.A(net1310),
    .B(_01119_),
    .X(_01125_));
 sky130_fd_sc_hd__a22o_1 _05150_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[31] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1476),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_2 _05151_ (.A(net1310),
    .B(_01121_),
    .X(_01126_));
 sky130_fd_sc_hd__a21o_1 _05152_ (.A1(net1476),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.hware_req ),
    .X(_00083_));
 sky130_fd_sc_hd__a22o_1 _05153_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[30] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1483),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05154_ (.A1(net1483),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.hware_req ),
    .X(_00082_));
 sky130_fd_sc_hd__a22o_1 _05155_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[29] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1499),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05156_ (.A1(net1499),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.hware_req ),
    .X(_00080_));
 sky130_fd_sc_hd__a22o_1 _05157_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[28] ),
    .A2(net1839),
    .B1(_01125_),
    .B2(net1507),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05158_ (.A1(net1507),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.hware_req ),
    .X(_00079_));
 sky130_fd_sc_hd__a22o_1 _05159_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[27] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1514),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05160_ (.A1(net1512),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.hware_req ),
    .X(_00078_));
 sky130_fd_sc_hd__a22o_1 _05161_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[26] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1521),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05162_ (.A1(net1521),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.hware_req ),
    .X(_00077_));
 sky130_fd_sc_hd__a22o_1 _05163_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[25] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1528),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05164_ (.A1(net1528),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.hware_req ),
    .X(_00076_));
 sky130_fd_sc_hd__a22o_1 _05165_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[24] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.data_out ),
    .B1(_01125_),
    .B2(net1536),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05166_ (.A1(net1536),
    .A2(_01126_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.hware_req ),
    .X(_00075_));
 sky130_fd_sc_hd__and2_2 _05167_ (.A(net1316),
    .B(_01119_),
    .X(_01127_));
 sky130_fd_sc_hd__a22o_1 _05168_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[23] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1542),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__and2_2 _05169_ (.A(net1316),
    .B(_01121_),
    .X(_01128_));
 sky130_fd_sc_hd__a21o_1 _05170_ (.A1(net1542),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.hware_req ),
    .X(_00074_));
 sky130_fd_sc_hd__a22o_1 _05171_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[22] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1552),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05172_ (.A1(net1550),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.hware_req ),
    .X(_00073_));
 sky130_fd_sc_hd__a22o_1 _05173_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[21] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1559),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05174_ (.A1(net1559),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.hware_req ),
    .X(_00072_));
 sky130_fd_sc_hd__a22o_1 _05175_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[20] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1566),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05176_ (.A1(net1567),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.hware_req ),
    .X(_00071_));
 sky130_fd_sc_hd__a22o_1 _05177_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[19] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1581),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05178_ (.A1(net1581),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.hware_req ),
    .X(_00069_));
 sky130_fd_sc_hd__a22o_1 _05179_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[18] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1589),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05180_ (.A1(net1589),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.hware_req ),
    .X(_00068_));
 sky130_fd_sc_hd__a22o_1 _05181_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[17] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1598),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05182_ (.A1(net1599),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.hware_req ),
    .X(_00067_));
 sky130_fd_sc_hd__a22o_1 _05183_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[16] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.data_out ),
    .B1(_01127_),
    .B2(net1606),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05184_ (.A1(net1606),
    .A2(_01128_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.hware_req ),
    .X(_00066_));
 sky130_fd_sc_hd__a22o_1 _05185_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[15] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1614),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05186_ (.A1(net1614),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.hware_req ),
    .X(_00065_));
 sky130_fd_sc_hd__a22o_1 _05187_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[14] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1621),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05188_ (.A1(net1622),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.hware_req ),
    .X(_00064_));
 sky130_fd_sc_hd__a22o_1 _05189_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[13] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1629),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05190_ (.A1(net1629),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.hware_req ),
    .X(_00063_));
 sky130_fd_sc_hd__a22o_1 _05191_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[12] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1636),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05192_ (.A1(net1637),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.hware_req ),
    .X(_00062_));
 sky130_fd_sc_hd__a22o_1 _05193_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[11] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1643),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05194_ (.A1(net1643),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.hware_req ),
    .X(_00061_));
 sky130_fd_sc_hd__a22o_1 _05195_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[10] ),
    .A2(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.data_out ),
    .B1(_01120_),
    .B2(net1287),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05196_ (.A1(net1287),
    .A2(_01122_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.hware_req ),
    .X(_00060_));
 sky130_fd_sc_hd__nor2_2 _05197_ (.A(net1345),
    .B(net1346),
    .Y(_01129_));
 sky130_fd_sc_hd__or2_2 _05198_ (.A(net1345),
    .B(net1346),
    .X(_01130_));
 sky130_fd_sc_hd__nor2_2 _05199_ (.A(_00999_),
    .B(_01130_),
    .Y(_01131_));
 sky130_fd_sc_hd__and3_4 _05200_ (.A(net1254),
    .B(net1179),
    .C(net1214),
    .X(_01132_));
 sky130_fd_sc_hd__a31o_1 _05201_ (.A1(net1308),
    .A2(net1166),
    .A3(net698),
    .B1(net1201),
    .X(_00126_));
 sky130_fd_sc_hd__a31o_1 _05202_ (.A1(net1316),
    .A2(net1169),
    .A3(net700),
    .B1(net1203),
    .X(_00125_));
 sky130_fd_sc_hd__a31o_1 _05203_ (.A1(net1323),
    .A2(net1169),
    .A3(net700),
    .B1(net1203),
    .X(_00124_));
 sky130_fd_sc_hd__a31o_1 _05204_ (.A1(net1331),
    .A2(net1166),
    .A3(net698),
    .B1(net1201),
    .X(_00123_));
 sky130_fd_sc_hd__nor2_1 _05205_ (.A(_01115_),
    .B(_01130_),
    .Y(_01133_));
 sky130_fd_sc_hd__and3_1 _05206_ (.A(net1254),
    .B(net1161),
    .C(net1214),
    .X(_01134_));
 sky130_fd_sc_hd__a31o_1 _05207_ (.A1(net1308),
    .A2(net1166),
    .A3(net685),
    .B1(_00795_),
    .X(_00150_));
 sky130_fd_sc_hd__a31o_1 _05208_ (.A1(net1316),
    .A2(net1170),
    .A3(net687),
    .B1(_00795_),
    .X(_00149_));
 sky130_fd_sc_hd__a31o_1 _05209_ (.A1(net1324),
    .A2(net1170),
    .A3(net687),
    .B1(_00795_),
    .X(_00148_));
 sky130_fd_sc_hd__a31o_1 _05210_ (.A1(net1331),
    .A2(net1167),
    .A3(net685),
    .B1(_00795_),
    .X(_00147_));
 sky130_fd_sc_hd__or2_1 _05211_ (.A(\u_glbl_reg.u_rtcclk.high_count[0] ),
    .B(\u_glbl_reg.u_rtcclk.high_count[1] ),
    .X(_01135_));
 sky130_fd_sc_hd__or2_1 _05212_ (.A(\u_glbl_reg.u_rtcclk.high_count[2] ),
    .B(_01135_),
    .X(_01136_));
 sky130_fd_sc_hd__or2_1 _05213_ (.A(\u_glbl_reg.u_rtcclk.high_count[3] ),
    .B(_01136_),
    .X(_01137_));
 sky130_fd_sc_hd__nor2_2 _05214_ (.A(\u_glbl_reg.u_rtcclk.high_count[4] ),
    .B(_01137_),
    .Y(_00194_));
 sky130_fd_sc_hd__nor2_1 _05215_ (.A(\u_glbl_reg.u_rtcclk.low_count[1] ),
    .B(\u_glbl_reg.u_rtcclk.low_count[0] ),
    .Y(_01138_));
 sky130_fd_sc_hd__or3_1 _05216_ (.A(\u_glbl_reg.u_rtcclk.low_count[1] ),
    .B(\u_glbl_reg.u_rtcclk.low_count[0] ),
    .C(\u_glbl_reg.u_rtcclk.low_count[2] ),
    .X(_01139_));
 sky130_fd_sc_hd__or2_1 _05217_ (.A(\u_glbl_reg.u_rtcclk.low_count[3] ),
    .B(_01139_),
    .X(_01140_));
 sky130_fd_sc_hd__inv_2 _05218_ (.A(_01140_),
    .Y(_01141_));
 sky130_fd_sc_hd__nor2_1 _05219_ (.A(\u_glbl_reg.u_rtcclk.low_count[4] ),
    .B(_01140_),
    .Y(_01142_));
 sky130_fd_sc_hd__or2_2 _05220_ (.A(\u_glbl_reg.u_rtcclk.low_count[4] ),
    .B(_01140_),
    .X(_01143_));
 sky130_fd_sc_hd__nand2_1 _05221_ (.A(_00194_),
    .B(_01143_),
    .Y(_00193_));
 sky130_fd_sc_hd__and2_4 _05222_ (.A(net1345),
    .B(net1346),
    .X(_01144_));
 sky130_fd_sc_hd__nand2_8 _05223_ (.A(net1255),
    .B(_01144_),
    .Y(_01145_));
 sky130_fd_sc_hd__nor2_8 _05224_ (.A(_00999_),
    .B(_01145_),
    .Y(_01146_));
 sky130_fd_sc_hd__a311o_1 _05225_ (.A1(net1308),
    .A2(net1166),
    .A3(net681),
    .B1(_00795_),
    .C1(_00796_),
    .X(_00236_));
 sky130_fd_sc_hd__and3_2 _05226_ (.A(net775),
    .B(net1170),
    .C(net683),
    .X(_01147_));
 sky130_fd_sc_hd__a21o_1 _05227_ (.A1(net1308),
    .A2(_01147_),
    .B1(_00796_),
    .X(_00235_));
 sky130_fd_sc_hd__a21o_1 _05228_ (.A1(net1316),
    .A2(_01147_),
    .B1(_00796_),
    .X(_00234_));
 sky130_fd_sc_hd__a21o_1 _05229_ (.A1(net1324),
    .A2(_01147_),
    .B1(_00796_),
    .X(_00233_));
 sky130_fd_sc_hd__a21o_1 _05230_ (.A1(net1331),
    .A2(_01147_),
    .B1(_00796_),
    .X(_00232_));
 sky130_fd_sc_hd__or2_1 _05231_ (.A(\u_glbl_reg.u_usbclk.high_count[0] ),
    .B(\u_glbl_reg.u_usbclk.high_count[1] ),
    .X(_01148_));
 sky130_fd_sc_hd__or2_1 _05232_ (.A(\u_glbl_reg.u_usbclk.high_count[2] ),
    .B(_01148_),
    .X(_01149_));
 sky130_fd_sc_hd__or2_1 _05233_ (.A(\u_glbl_reg.u_usbclk.high_count[3] ),
    .B(_01149_),
    .X(_01150_));
 sky130_fd_sc_hd__nor2_2 _05234_ (.A(\u_glbl_reg.u_usbclk.high_count[4] ),
    .B(_01150_),
    .Y(_00244_));
 sky130_fd_sc_hd__nor2_1 _05235_ (.A(\u_glbl_reg.u_usbclk.low_count[1] ),
    .B(\u_glbl_reg.u_usbclk.low_count[0] ),
    .Y(_01151_));
 sky130_fd_sc_hd__or3_1 _05236_ (.A(\u_glbl_reg.u_usbclk.low_count[1] ),
    .B(\u_glbl_reg.u_usbclk.low_count[0] ),
    .C(\u_glbl_reg.u_usbclk.low_count[2] ),
    .X(_01152_));
 sky130_fd_sc_hd__or2_1 _05237_ (.A(\u_glbl_reg.u_usbclk.low_count[3] ),
    .B(_01152_),
    .X(_01153_));
 sky130_fd_sc_hd__inv_2 _05238_ (.A(_01153_),
    .Y(_01154_));
 sky130_fd_sc_hd__nor2_1 _05239_ (.A(\u_glbl_reg.u_usbclk.low_count[4] ),
    .B(_01153_),
    .Y(_01155_));
 sky130_fd_sc_hd__or2_2 _05240_ (.A(\u_glbl_reg.u_usbclk.low_count[4] ),
    .B(_01153_),
    .X(_01156_));
 sky130_fd_sc_hd__nand2_1 _05241_ (.A(_00244_),
    .B(_01156_),
    .Y(_00243_));
 sky130_fd_sc_hd__nand2_1 _05242_ (.A(_00807_),
    .B(\u_ws281x.cfg_reset_period[5] ),
    .Y(_01157_));
 sky130_fd_sc_hd__a22o_1 _05243_ (.A1(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .A2(_00814_),
    .B1(_00821_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .X(_01158_));
 sky130_fd_sc_hd__a221o_1 _05244_ (.A1(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .A2(_00818_),
    .B1(_00819_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .C1(_01158_),
    .X(_01159_));
 sky130_fd_sc_hd__o22ai_1 _05245_ (.A1(_00805_),
    .A2(\u_ws281x.cfg_reset_period[4] ),
    .B1(_00821_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .Y(_01160_));
 sky130_fd_sc_hd__a221o_1 _05246_ (.A1(_00802_),
    .A2(\u_ws281x.cfg_reset_period[2] ),
    .B1(\u_ws281x.cfg_reset_period[4] ),
    .B2(_00805_),
    .C1(_01160_),
    .X(_01161_));
 sky130_fd_sc_hd__nor2_1 _05247_ (.A(_01159_),
    .B(_01161_),
    .Y(_01162_));
 sky130_fd_sc_hd__o2bb2a_1 _05248_ (.A1_N(\u_ws281x.u_txd_0.clk_cnt[12] ),
    .A2_N(_00822_),
    .B1(_00814_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .X(_01163_));
 sky130_fd_sc_hd__xnor2_1 _05249_ (.A(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .B(\u_ws281x.cfg_reset_period[10] ),
    .Y(_01164_));
 sky130_fd_sc_hd__o221a_1 _05250_ (.A1(_00802_),
    .A2(\u_ws281x.cfg_reset_period[2] ),
    .B1(_00823_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .C1(_01164_),
    .X(_01165_));
 sky130_fd_sc_hd__o221a_1 _05251_ (.A1(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .A2(_00818_),
    .B1(_00819_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .C1(_01163_),
    .X(_01166_));
 sky130_fd_sc_hd__xnor2_1 _05252_ (.A(\u_ws281x.u_txd_0.clk_cnt[14] ),
    .B(\u_ws281x.cfg_reset_period[14] ),
    .Y(_01167_));
 sky130_fd_sc_hd__o221a_1 _05253_ (.A1(_00808_),
    .A2(\u_ws281x.cfg_reset_period[6] ),
    .B1(\u_ws281x.cfg_reset_period[9] ),
    .B2(_00812_),
    .C1(_01167_),
    .X(_01168_));
 sky130_fd_sc_hd__a22o_1 _05254_ (.A1(_00808_),
    .A2(\u_ws281x.cfg_reset_period[6] ),
    .B1(_00824_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[15] ),
    .X(_01169_));
 sky130_fd_sc_hd__a22o_1 _05255_ (.A1(_00798_),
    .A2(\u_ws281x.cfg_reset_period[0] ),
    .B1(\u_ws281x.cfg_reset_period[3] ),
    .B2(_00804_),
    .X(_01170_));
 sky130_fd_sc_hd__a211oi_1 _05256_ (.A1(\u_ws281x.u_txd_0.clk_cnt[5] ),
    .A2(_00816_),
    .B1(_01169_),
    .C1(_01170_),
    .Y(_01171_));
 sky130_fd_sc_hd__o2bb2a_1 _05257_ (.A1_N(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .A2_N(_00823_),
    .B1(_00820_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .X(_01172_));
 sky130_fd_sc_hd__o221a_1 _05258_ (.A1(\u_ws281x.u_txd_0.clk_cnt[12] ),
    .A2(_00822_),
    .B1(_00824_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[15] ),
    .C1(_01157_),
    .X(_01173_));
 sky130_fd_sc_hd__o2111a_1 _05259_ (.A1(_00804_),
    .A2(\u_ws281x.cfg_reset_period[3] ),
    .B1(_01171_),
    .C1(_01172_),
    .D1(_01173_),
    .X(_01174_));
 sky130_fd_sc_hd__o211a_1 _05260_ (.A1(_00798_),
    .A2(\u_ws281x.cfg_reset_period[0] ),
    .B1(_01168_),
    .C1(_01174_),
    .X(_01175_));
 sky130_fd_sc_hd__and4_1 _05261_ (.A(_01162_),
    .B(_01165_),
    .C(_01166_),
    .D(_01175_),
    .X(_01176_));
 sky130_fd_sc_hd__inv_2 _05262_ (.A(_01176_),
    .Y(_01177_));
 sky130_fd_sc_hd__and2_1 _05263_ (.A(\u_ws281x.port0_enb ),
    .B(_01176_),
    .X(_01178_));
 sky130_fd_sc_hd__nor2_1 _05264_ (.A(\u_ws281x.u_txd_0.state ),
    .B(_01178_),
    .Y(_01179_));
 sky130_fd_sc_hd__a22o_1 _05265_ (.A1(\u_ws281x.cfg_clk_period[5] ),
    .A2(_00807_),
    .B1(_00811_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .X(_01180_));
 sky130_fd_sc_hd__a2bb2o_1 _05266_ (.A1_N(\u_ws281x.cfg_clk_period[4] ),
    .A2_N(_00805_),
    .B1(\u_ws281x.cfg_clk_period[3] ),
    .B2(_00804_),
    .X(_01181_));
 sky130_fd_sc_hd__or4_1 _05267_ (.A(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[12] ),
    .C(\u_ws281x.u_txd_0.clk_cnt[15] ),
    .D(\u_ws281x.u_txd_0.clk_cnt[14] ),
    .X(_01182_));
 sky130_fd_sc_hd__a211o_1 _05268_ (.A1(_00806_),
    .A2(\u_ws281x.u_txd_0.clk_cnt[5] ),
    .B1(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .C1(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .X(_01183_));
 sky130_fd_sc_hd__or4_1 _05269_ (.A(_01180_),
    .B(_01181_),
    .C(_01182_),
    .D(_01183_),
    .X(_01184_));
 sky130_fd_sc_hd__a22o_1 _05270_ (.A1(_00799_),
    .A2(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .B1(\u_ws281x.cfg_clk_period[9] ),
    .B2(_00812_),
    .X(_01185_));
 sky130_fd_sc_hd__a221o_1 _05271_ (.A1(_00801_),
    .A2(\u_ws281x.u_txd_0.clk_cnt[2] ),
    .B1(\u_ws281x.cfg_clk_period[6] ),
    .B2(_00808_),
    .C1(_01185_),
    .X(_01186_));
 sky130_fd_sc_hd__a22o_1 _05272_ (.A1(_00797_),
    .A2(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .B1(\u_ws281x.cfg_clk_period[1] ),
    .B2(_00800_),
    .X(_01187_));
 sky130_fd_sc_hd__a221o_1 _05273_ (.A1(\u_ws281x.cfg_clk_period[4] ),
    .A2(_00805_),
    .B1(\u_ws281x.cfg_clk_period[8] ),
    .B2(_00810_),
    .C1(_01187_),
    .X(_01188_));
 sky130_fd_sc_hd__nor2_1 _05274_ (.A(\u_ws281x.cfg_clk_period[6] ),
    .B(_00808_),
    .Y(_01189_));
 sky130_fd_sc_hd__a221o_1 _05275_ (.A1(\u_ws281x.cfg_clk_period[0] ),
    .A2(_00798_),
    .B1(_00803_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[3] ),
    .C1(_01189_),
    .X(_01190_));
 sky130_fd_sc_hd__o2bb2a_1 _05276_ (.A1_N(_00809_),
    .A2_N(\u_ws281x.cfg_clk_period[7] ),
    .B1(\u_ws281x.u_txd_0.clk_cnt[2] ),
    .B2(_00801_),
    .X(_01191_));
 sky130_fd_sc_hd__o221a_1 _05277_ (.A1(\u_ws281x.cfg_clk_period[7] ),
    .A2(_00809_),
    .B1(\u_ws281x.cfg_clk_period[8] ),
    .B2(_00810_),
    .C1(_01191_),
    .X(_01192_));
 sky130_fd_sc_hd__or4b_1 _05278_ (.A(_01186_),
    .B(_01188_),
    .C(_01190_),
    .D_N(_01192_),
    .X(_01193_));
 sky130_fd_sc_hd__or2_1 _05279_ (.A(_01184_),
    .B(_01193_),
    .X(_01194_));
 sky130_fd_sc_hd__nand2_1 _05280_ (.A(\u_ws281x.u_txd_0.state ),
    .B(_01194_),
    .Y(_01195_));
 sky130_fd_sc_hd__inv_2 _05281_ (.A(_01195_),
    .Y(_01196_));
 sky130_fd_sc_hd__or3_2 _05282_ (.A(\u_ws281x.u_txd_0.bit_cnt[0] ),
    .B(\u_ws281x.u_txd_0.bit_cnt[1] ),
    .C(\u_ws281x.u_txd_0.bit_cnt[2] ),
    .X(_01197_));
 sky130_fd_sc_hd__o31ai_4 _05283_ (.A1(\u_ws281x.u_txd_0.bit_cnt[3] ),
    .A2(\u_ws281x.u_txd_0.bit_cnt[4] ),
    .A3(_01197_),
    .B1(net2099),
    .Y(_01198_));
 sky130_fd_sc_hd__inv_2 _05284_ (.A(net574),
    .Y(_01199_));
 sky130_fd_sc_hd__o211ai_1 _05285_ (.A1(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .A2(_01179_),
    .B1(_01195_),
    .C1(net574),
    .Y(_04681_));
 sky130_fd_sc_hd__xor2_1 _05286_ (.A(\u_ws281x.cfg_reset_period[10] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[10] ),
    .X(_01200_));
 sky130_fd_sc_hd__a221o_1 _05287_ (.A1(\u_ws281x.cfg_reset_period[2] ),
    .A2(_00828_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[13] ),
    .B2(_00823_),
    .C1(_01200_),
    .X(_01201_));
 sky130_fd_sc_hd__o22a_1 _05288_ (.A1(\u_ws281x.cfg_reset_period[1] ),
    .A2(_00827_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .B2(_00822_),
    .X(_01202_));
 sky130_fd_sc_hd__a22o_1 _05289_ (.A1(\u_ws281x.cfg_reset_period[4] ),
    .A2(_00830_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[11] ),
    .B2(_00821_),
    .X(_01203_));
 sky130_fd_sc_hd__o22a_1 _05290_ (.A1(\u_ws281x.cfg_reset_period[2] ),
    .A2(_00828_),
    .B1(_00830_),
    .B2(\u_ws281x.cfg_reset_period[4] ),
    .X(_01204_));
 sky130_fd_sc_hd__o22a_1 _05291_ (.A1(_00814_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[11] ),
    .B2(_00821_),
    .X(_01205_));
 sky130_fd_sc_hd__o221a_1 _05292_ (.A1(\u_ws281x.cfg_reset_period[7] ),
    .A2(_00833_),
    .B1(_00834_),
    .B2(\u_ws281x.cfg_reset_period[8] ),
    .C1(_01202_),
    .X(_01206_));
 sky130_fd_sc_hd__o221a_1 _05293_ (.A1(_00818_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[8] ),
    .B2(_00819_),
    .C1(_01205_),
    .X(_01207_));
 sky130_fd_sc_hd__and4bb_1 _05294_ (.A_N(_01201_),
    .B_N(_01203_),
    .C(_01204_),
    .D(_01207_),
    .X(_01208_));
 sky130_fd_sc_hd__xnor2_1 _05295_ (.A(\u_ws281x.cfg_reset_period[14] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[14] ),
    .Y(_01209_));
 sky130_fd_sc_hd__o221a_1 _05296_ (.A1(_00817_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[6] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .B2(_00820_),
    .C1(_01209_),
    .X(_01210_));
 sky130_fd_sc_hd__o22a_1 _05297_ (.A1(\u_ws281x.cfg_reset_period[6] ),
    .A2(_00832_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[15] ),
    .B2(_00824_),
    .X(_01211_));
 sky130_fd_sc_hd__o22a_1 _05298_ (.A1(\u_ws281x.cfg_reset_period[9] ),
    .A2(_00835_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[13] ),
    .B2(_00823_),
    .X(_01212_));
 sky130_fd_sc_hd__a22o_1 _05299_ (.A1(_00822_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[15] ),
    .B2(_00824_),
    .X(_01213_));
 sky130_fd_sc_hd__a221o_1 _05300_ (.A1(\u_ws281x.cfg_reset_period[0] ),
    .A2(_00826_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .B2(_00816_),
    .C1(_01213_),
    .X(_01214_));
 sky130_fd_sc_hd__o221a_1 _05301_ (.A1(\u_ws281x.cfg_reset_period[3] ),
    .A2(_00829_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .B2(_00816_),
    .C1(_01211_),
    .X(_01215_));
 sky130_fd_sc_hd__o221a_1 _05302_ (.A1(\u_ws281x.cfg_reset_period[0] ),
    .A2(_00826_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .B2(_00815_),
    .C1(_01212_),
    .X(_01216_));
 sky130_fd_sc_hd__and3_1 _05303_ (.A(_01210_),
    .B(_01215_),
    .C(_01216_),
    .X(_01217_));
 sky130_fd_sc_hd__and2b_1 _05304_ (.A_N(_01214_),
    .B(_01217_),
    .X(_01218_));
 sky130_fd_sc_hd__and3_1 _05305_ (.A(_01206_),
    .B(_01208_),
    .C(_01218_),
    .X(_01219_));
 sky130_fd_sc_hd__and2_1 _05306_ (.A(\u_ws281x.port1_enb ),
    .B(_01219_),
    .X(_01220_));
 sky130_fd_sc_hd__nor2_1 _05307_ (.A(\u_ws281x.u_txd_1.state ),
    .B(_01220_),
    .Y(_01221_));
 sky130_fd_sc_hd__nor2_1 _05308_ (.A(\u_ws281x.cfg_clk_period[8] ),
    .B(_00834_),
    .Y(_01222_));
 sky130_fd_sc_hd__or4_1 _05309_ (.A(\u_ws281x.u_txd_1.clk_cnt[13] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .C(\u_ws281x.u_txd_1.clk_cnt[15] ),
    .D(\u_ws281x.u_txd_1.clk_cnt[14] ),
    .X(_01223_));
 sky130_fd_sc_hd__a22o_1 _05310_ (.A1(\u_ws281x.cfg_clk_period[1] ),
    .A2(_00827_),
    .B1(_00835_),
    .B2(\u_ws281x.cfg_clk_period[9] ),
    .X(_01224_));
 sky130_fd_sc_hd__a2bb2o_1 _05311_ (.A1_N(_00832_),
    .A2_N(\u_ws281x.cfg_clk_period[6] ),
    .B1(_00801_),
    .B2(\u_ws281x.u_txd_1.clk_cnt[2] ),
    .X(_01225_));
 sky130_fd_sc_hd__xor2_1 _05312_ (.A(\u_ws281x.cfg_clk_period[4] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[4] ),
    .X(_01226_));
 sky130_fd_sc_hd__xor2_1 _05313_ (.A(\u_ws281x.cfg_clk_period[7] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .X(_01227_));
 sky130_fd_sc_hd__xor2_1 _05314_ (.A(\u_ws281x.cfg_clk_period[5] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .X(_01228_));
 sky130_fd_sc_hd__or4_1 _05315_ (.A(_01223_),
    .B(_01226_),
    .C(_01227_),
    .D(_01228_),
    .X(_01229_));
 sky130_fd_sc_hd__a22o_1 _05316_ (.A1(\u_ws281x.cfg_clk_period[2] ),
    .A2(_00828_),
    .B1(_00829_),
    .B2(\u_ws281x.cfg_clk_period[3] ),
    .X(_01230_));
 sky130_fd_sc_hd__a211o_1 _05317_ (.A1(_00799_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[11] ),
    .C1(\u_ws281x.u_txd_1.clk_cnt[10] ),
    .X(_01231_));
 sky130_fd_sc_hd__a221o_1 _05318_ (.A1(\u_ws281x.cfg_clk_period[0] ),
    .A2(_00826_),
    .B1(_00832_),
    .B2(\u_ws281x.cfg_clk_period[6] ),
    .C1(_01222_),
    .X(_01232_));
 sky130_fd_sc_hd__a221o_1 _05319_ (.A1(_00797_),
    .A2(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .B2(_00803_),
    .C1(_01232_),
    .X(_01233_));
 sky130_fd_sc_hd__a221o_1 _05320_ (.A1(\u_ws281x.cfg_clk_period[8] ),
    .A2(_00834_),
    .B1(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .B2(_00811_),
    .C1(_01233_),
    .X(_01234_));
 sky130_fd_sc_hd__or4_1 _05321_ (.A(_01224_),
    .B(_01225_),
    .C(_01229_),
    .D(_01234_),
    .X(_01235_));
 sky130_fd_sc_hd__or3_2 _05322_ (.A(_01230_),
    .B(_01231_),
    .C(_01235_),
    .X(_01236_));
 sky130_fd_sc_hd__nand2_1 _05323_ (.A(\u_ws281x.u_txd_1.state ),
    .B(_01236_),
    .Y(_01237_));
 sky130_fd_sc_hd__or3_2 _05324_ (.A(\u_ws281x.u_txd_1.bit_cnt[0] ),
    .B(\u_ws281x.u_txd_1.bit_cnt[1] ),
    .C(\u_ws281x.u_txd_1.bit_cnt[2] ),
    .X(_01238_));
 sky130_fd_sc_hd__o31ai_4 _05325_ (.A1(\u_ws281x.u_txd_1.bit_cnt[3] ),
    .A2(\u_ws281x.u_txd_1.bit_cnt[4] ),
    .A3(_01238_),
    .B1(net2089),
    .Y(_01239_));
 sky130_fd_sc_hd__inv_2 _05326_ (.A(net570),
    .Y(_01240_));
 sky130_fd_sc_hd__o211ai_1 _05327_ (.A1(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .A2(_01221_),
    .B1(_01237_),
    .C1(net570),
    .Y(_04687_));
 sky130_fd_sc_hd__a22o_1 _05328_ (.A1(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ),
    .A2(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.data_out ),
    .B1(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ),
    .B2(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[1].u_bit_reg.data_out ),
    .X(_01241_));
 sky130_fd_sc_hd__a221o_4 _05329_ (.A1(net2168),
    .A2(net1834),
    .B1(_01123_),
    .B2(net1450),
    .C1(_01241_),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05330_ (.A1(net1452),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ),
    .X(_00086_));
 sky130_fd_sc_hd__a31o_1 _05331_ (.A1(net1332),
    .A2(net1458),
    .A3(_01119_),
    .B1(\u_glbl_reg.usb_intr_ss ),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05332_ (.A1(net1461),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.hware_req ),
    .X(_00085_));
 sky130_fd_sc_hd__a31o_1 _05333_ (.A1(net1332),
    .A2(net1467),
    .A3(_01119_),
    .B1(\u_glbl_reg.i2cm_intr_ss ),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05334_ (.A1(net1467),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.hware_req ),
    .X(_00084_));
 sky130_fd_sc_hd__or3_1 _05335_ (.A(\u_timer.u_timer_2.timer_counter[0] ),
    .B(\u_timer.u_timer_2.timer_counter[1] ),
    .C(\u_timer.u_timer_2.timer_counter[2] ),
    .X(_01242_));
 sky130_fd_sc_hd__or2_1 _05336_ (.A(\u_timer.u_timer_2.timer_counter[3] ),
    .B(_01242_),
    .X(_01243_));
 sky130_fd_sc_hd__or3_1 _05337_ (.A(\u_timer.u_timer_2.timer_counter[5] ),
    .B(\u_timer.u_timer_2.timer_counter[4] ),
    .C(_01243_),
    .X(_01244_));
 sky130_fd_sc_hd__or2_1 _05338_ (.A(\u_timer.u_timer_2.timer_counter[6] ),
    .B(_01244_),
    .X(_01245_));
 sky130_fd_sc_hd__or3_1 _05339_ (.A(\u_timer.u_timer_2.timer_counter[7] ),
    .B(\u_timer.u_timer_2.timer_counter[8] ),
    .C(_01245_),
    .X(_01246_));
 sky130_fd_sc_hd__or2_1 _05340_ (.A(\u_timer.u_timer_2.timer_counter[9] ),
    .B(_01246_),
    .X(_01247_));
 sky130_fd_sc_hd__or3_1 _05341_ (.A(\u_timer.u_timer_2.timer_counter[11] ),
    .B(\u_timer.u_timer_2.timer_counter[10] ),
    .C(_01247_),
    .X(_01248_));
 sky130_fd_sc_hd__or2_1 _05342_ (.A(\u_timer.u_timer_2.timer_counter[12] ),
    .B(_01248_),
    .X(_01249_));
 sky130_fd_sc_hd__or3_1 _05343_ (.A(\u_timer.u_timer_2.timer_counter[13] ),
    .B(\u_timer.u_timer_2.timer_counter[14] ),
    .C(_01249_),
    .X(_01250_));
 sky130_fd_sc_hd__nor2_1 _05344_ (.A(\u_timer.u_timer_2.timer_counter[15] ),
    .B(_01250_),
    .Y(\u_timer.u_timer_2.timer_hit ));
 sky130_fd_sc_hd__a32o_2 _05345_ (.A1(_00841_),
    .A2(\u_timer.cfg_timer2[16] ),
    .A3(\u_timer.u_timer_2.timer_hit ),
    .B1(_01123_),
    .B2(net1494),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05346_ (.A1(net1494),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .X(_00081_));
 sky130_fd_sc_hd__or3_1 _05347_ (.A(\u_timer.u_timer_1.timer_counter[0] ),
    .B(\u_timer.u_timer_1.timer_counter[1] ),
    .C(\u_timer.u_timer_1.timer_counter[2] ),
    .X(_01251_));
 sky130_fd_sc_hd__or2_1 _05348_ (.A(\u_timer.u_timer_1.timer_counter[3] ),
    .B(_01251_),
    .X(_01252_));
 sky130_fd_sc_hd__or3_1 _05349_ (.A(\u_timer.u_timer_1.timer_counter[5] ),
    .B(\u_timer.u_timer_1.timer_counter[4] ),
    .C(_01252_),
    .X(_01253_));
 sky130_fd_sc_hd__or2_1 _05350_ (.A(\u_timer.u_timer_1.timer_counter[6] ),
    .B(_01253_),
    .X(_01254_));
 sky130_fd_sc_hd__or3_1 _05351_ (.A(\u_timer.u_timer_1.timer_counter[7] ),
    .B(\u_timer.u_timer_1.timer_counter[8] ),
    .C(_01254_),
    .X(_01255_));
 sky130_fd_sc_hd__or2_1 _05352_ (.A(\u_timer.u_timer_1.timer_counter[9] ),
    .B(_01255_),
    .X(_01256_));
 sky130_fd_sc_hd__or3_1 _05353_ (.A(\u_timer.u_timer_1.timer_counter[11] ),
    .B(\u_timer.u_timer_1.timer_counter[10] ),
    .C(_01256_),
    .X(_01257_));
 sky130_fd_sc_hd__or2_1 _05354_ (.A(\u_timer.u_timer_1.timer_counter[12] ),
    .B(_01257_),
    .X(_01258_));
 sky130_fd_sc_hd__or3_1 _05355_ (.A(\u_timer.u_timer_1.timer_counter[13] ),
    .B(\u_timer.u_timer_1.timer_counter[14] ),
    .C(_01258_),
    .X(_01259_));
 sky130_fd_sc_hd__nor2_1 _05356_ (.A(\u_timer.u_timer_1.timer_counter[15] ),
    .B(_01259_),
    .Y(\u_timer.u_timer_1.timer_hit ));
 sky130_fd_sc_hd__a32o_2 _05357_ (.A1(_00844_),
    .A2(\u_timer.cfg_timer1[16] ),
    .A3(\u_timer.u_timer_1.timer_hit ),
    .B1(_01123_),
    .B2(net1577),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05358_ (.A1(net1577),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .X(_00070_));
 sky130_fd_sc_hd__or3_1 _05359_ (.A(\u_timer.u_timer_0.timer_counter[0] ),
    .B(\u_timer.u_timer_0.timer_counter[1] ),
    .C(\u_timer.u_timer_0.timer_counter[2] ),
    .X(_01260_));
 sky130_fd_sc_hd__or2_1 _05360_ (.A(\u_timer.u_timer_0.timer_counter[3] ),
    .B(_01260_),
    .X(_01261_));
 sky130_fd_sc_hd__or3_1 _05361_ (.A(\u_timer.u_timer_0.timer_counter[5] ),
    .B(\u_timer.u_timer_0.timer_counter[4] ),
    .C(_01261_),
    .X(_01262_));
 sky130_fd_sc_hd__or2_1 _05362_ (.A(\u_timer.u_timer_0.timer_counter[6] ),
    .B(_01262_),
    .X(_01263_));
 sky130_fd_sc_hd__or3_1 _05363_ (.A(\u_timer.u_timer_0.timer_counter[7] ),
    .B(\u_timer.u_timer_0.timer_counter[8] ),
    .C(_01263_),
    .X(_01264_));
 sky130_fd_sc_hd__or2_1 _05364_ (.A(\u_timer.u_timer_0.timer_counter[9] ),
    .B(_01264_),
    .X(_01265_));
 sky130_fd_sc_hd__or3_1 _05365_ (.A(\u_timer.u_timer_0.timer_counter[11] ),
    .B(\u_timer.u_timer_0.timer_counter[10] ),
    .C(_01265_),
    .X(_01266_));
 sky130_fd_sc_hd__or2_1 _05366_ (.A(\u_timer.u_timer_0.timer_counter[12] ),
    .B(_01266_),
    .X(_01267_));
 sky130_fd_sc_hd__or3_1 _05367_ (.A(\u_timer.u_timer_0.timer_counter[13] ),
    .B(\u_timer.u_timer_0.timer_counter[14] ),
    .C(_01267_),
    .X(_01268_));
 sky130_fd_sc_hd__nor2_1 _05368_ (.A(\u_timer.u_timer_0.timer_counter[15] ),
    .B(_01268_),
    .Y(\u_timer.u_timer_0.timer_hit ));
 sky130_fd_sc_hd__a32o_2 _05369_ (.A1(_00847_),
    .A2(\u_timer.cfg_timer0[16] ),
    .A3(\u_timer.u_timer_0.timer_hit ),
    .B1(_01123_),
    .B2(net1299),
    .X(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__a21o_1 _05370_ (.A1(net1298),
    .A2(_01124_),
    .B1(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .X(_00059_));
 sky130_fd_sc_hd__and3b_1 _05371_ (.A_N(net1374),
    .B(net1340),
    .C(net1342),
    .X(_01269_));
 sky130_fd_sc_hd__and3_2 _05372_ (.A(net1416),
    .B(_01002_),
    .C(_01269_),
    .X(_01270_));
 sky130_fd_sc_hd__and4_2 _05373_ (.A(\u_ws281x.reg_ack ),
    .B(_00850_),
    .C(net714),
    .D(_01270_),
    .X(_00589_));
 sky130_fd_sc_hd__xnor2_1 _05374_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.wr_ptr ),
    .B(net1084),
    .Y(_01271_));
 sky130_fd_sc_hd__nor3_1 _05375_ (.A(_00849_),
    .B(_00589_),
    .C(_01271_),
    .Y(_00587_));
 sky130_fd_sc_hd__and3_1 _05376_ (.A(_00849_),
    .B(_00589_),
    .C(_01271_),
    .X(_00588_));
 sky130_fd_sc_hd__or2_1 _05377_ (.A(_00587_),
    .B(_00588_),
    .X(_00591_));
 sky130_fd_sc_hd__and4_1 _05378_ (.A(\u_ws281x.reg_ack ),
    .B(_00852_),
    .C(net710),
    .D(_01270_),
    .X(_00582_));
 sky130_fd_sc_hd__xnor2_1 _05379_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.wr_ptr ),
    .B(net1080),
    .Y(_01272_));
 sky130_fd_sc_hd__nor3_1 _05380_ (.A(_00851_),
    .B(_00582_),
    .C(_01272_),
    .Y(_00580_));
 sky130_fd_sc_hd__and3_1 _05381_ (.A(_00851_),
    .B(_00582_),
    .C(_01272_),
    .X(_00581_));
 sky130_fd_sc_hd__or2_1 _05382_ (.A(_00580_),
    .B(_00581_),
    .X(_00584_));
 sky130_fd_sc_hd__o22a_1 _05383_ (.A1(\u_ws281x.u_txd_0.state ),
    .A2(_01178_),
    .B1(_01194_),
    .B2(net574),
    .X(_00649_));
 sky130_fd_sc_hd__or3b_1 _05384_ (.A(net734),
    .B(\u_ws281x.u_txd_0.state ),
    .C_N(_01178_),
    .X(_00650_));
 sky130_fd_sc_hd__or2_1 _05385_ (.A(_00805_),
    .B(\u_ws281x.cfg_th1_period[4] ),
    .X(_01273_));
 sky130_fd_sc_hd__nand2_1 _05386_ (.A(\u_ws281x.u_txd_0.clk_cnt[3] ),
    .B(_00854_),
    .Y(_01274_));
 sky130_fd_sc_hd__or2_1 _05387_ (.A(_00798_),
    .B(\u_ws281x.cfg_th1_period[0] ),
    .X(_01275_));
 sky130_fd_sc_hd__nor2_1 _05388_ (.A(_00812_),
    .B(\u_ws281x.cfg_th1_period[9] ),
    .Y(_01276_));
 sky130_fd_sc_hd__a221o_1 _05389_ (.A1(_00798_),
    .A2(\u_ws281x.cfg_th1_period[0] ),
    .B1(_00855_),
    .B2(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .C1(_01276_),
    .X(_01277_));
 sky130_fd_sc_hd__a22o_1 _05390_ (.A1(_00800_),
    .A2(\u_ws281x.cfg_th1_period[1] ),
    .B1(_01275_),
    .B2(_01277_),
    .X(_01278_));
 sky130_fd_sc_hd__o221a_1 _05391_ (.A1(_00800_),
    .A2(\u_ws281x.cfg_th1_period[1] ),
    .B1(\u_ws281x.cfg_th1_period[2] ),
    .B2(_00802_),
    .C1(_01278_),
    .X(_01279_));
 sky130_fd_sc_hd__a221o_1 _05392_ (.A1(_00804_),
    .A2(\u_ws281x.cfg_th1_period[3] ),
    .B1(\u_ws281x.cfg_th1_period[2] ),
    .B2(_00802_),
    .C1(_01279_),
    .X(_01280_));
 sky130_fd_sc_hd__a22o_1 _05393_ (.A1(_00805_),
    .A2(\u_ws281x.cfg_th1_period[4] ),
    .B1(_01274_),
    .B2(_01280_),
    .X(_01281_));
 sky130_fd_sc_hd__a22o_1 _05394_ (.A1(_00807_),
    .A2(\u_ws281x.cfg_th1_period[5] ),
    .B1(_01273_),
    .B2(_01281_),
    .X(_01282_));
 sky130_fd_sc_hd__o221a_1 _05395_ (.A1(_00808_),
    .A2(\u_ws281x.cfg_th1_period[6] ),
    .B1(\u_ws281x.cfg_th1_period[5] ),
    .B2(_00807_),
    .C1(_01282_),
    .X(_01283_));
 sky130_fd_sc_hd__a221o_1 _05396_ (.A1(_00809_),
    .A2(\u_ws281x.cfg_th1_period[7] ),
    .B1(\u_ws281x.cfg_th1_period[6] ),
    .B2(_00808_),
    .C1(_01283_),
    .X(_01284_));
 sky130_fd_sc_hd__o221a_1 _05397_ (.A1(_00809_),
    .A2(\u_ws281x.cfg_th1_period[7] ),
    .B1(\u_ws281x.cfg_th1_period[8] ),
    .B2(_00810_),
    .C1(_01284_),
    .X(_01285_));
 sky130_fd_sc_hd__a22o_1 _05398_ (.A1(_00812_),
    .A2(\u_ws281x.cfg_th1_period[9] ),
    .B1(\u_ws281x.cfg_th1_period[8] ),
    .B2(_00810_),
    .X(_01286_));
 sky130_fd_sc_hd__o21ba_1 _05399_ (.A1(_01285_),
    .A2(_01286_),
    .B1_N(_01276_),
    .X(_01287_));
 sky130_fd_sc_hd__o211a_1 _05400_ (.A1(_00798_),
    .A2(\u_ws281x.cfg_th0_period[0] ),
    .B1(_00853_),
    .C1(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .X(_01288_));
 sky130_fd_sc_hd__a221o_1 _05401_ (.A1(_00800_),
    .A2(\u_ws281x.cfg_th0_period[1] ),
    .B1(\u_ws281x.cfg_th0_period[0] ),
    .B2(_00798_),
    .C1(_01288_),
    .X(_01289_));
 sky130_fd_sc_hd__o221a_1 _05402_ (.A1(_00802_),
    .A2(\u_ws281x.cfg_th0_period[2] ),
    .B1(\u_ws281x.cfg_th0_period[1] ),
    .B2(_00800_),
    .C1(_01289_),
    .X(_01290_));
 sky130_fd_sc_hd__a221o_1 _05403_ (.A1(_00804_),
    .A2(\u_ws281x.cfg_th0_period[3] ),
    .B1(\u_ws281x.cfg_th0_period[2] ),
    .B2(_00802_),
    .C1(_01290_),
    .X(_01291_));
 sky130_fd_sc_hd__o221a_1 _05404_ (.A1(_00805_),
    .A2(\u_ws281x.cfg_th0_period[4] ),
    .B1(\u_ws281x.cfg_th0_period[3] ),
    .B2(_00804_),
    .C1(_01291_),
    .X(_01292_));
 sky130_fd_sc_hd__a221o_1 _05405_ (.A1(_00807_),
    .A2(\u_ws281x.cfg_th0_period[5] ),
    .B1(\u_ws281x.cfg_th0_period[4] ),
    .B2(_00805_),
    .C1(_01292_),
    .X(_01293_));
 sky130_fd_sc_hd__o221a_1 _05406_ (.A1(_00808_),
    .A2(\u_ws281x.cfg_th0_period[6] ),
    .B1(\u_ws281x.cfg_th0_period[5] ),
    .B2(_00807_),
    .C1(_01293_),
    .X(_01294_));
 sky130_fd_sc_hd__a221o_1 _05407_ (.A1(_00809_),
    .A2(\u_ws281x.cfg_th0_period[7] ),
    .B1(\u_ws281x.cfg_th0_period[6] ),
    .B2(_00808_),
    .C1(_01294_),
    .X(_01295_));
 sky130_fd_sc_hd__o221a_1 _05408_ (.A1(_00810_),
    .A2(\u_ws281x.cfg_th0_period[8] ),
    .B1(\u_ws281x.cfg_th0_period[7] ),
    .B2(_00809_),
    .C1(_01295_),
    .X(_01296_));
 sky130_fd_sc_hd__a221o_1 _05409_ (.A1(_00812_),
    .A2(\u_ws281x.cfg_th0_period[9] ),
    .B1(\u_ws281x.cfg_th0_period[8] ),
    .B2(_00810_),
    .C1(_01296_),
    .X(_01297_));
 sky130_fd_sc_hd__a21oi_1 _05410_ (.A1(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .A2(_00853_),
    .B1(\u_ws281x.u_txd_0.led_data[23] ),
    .Y(_01298_));
 sky130_fd_sc_hd__a22oi_2 _05411_ (.A1(\u_ws281x.u_txd_0.led_data[23] ),
    .A2(_01287_),
    .B1(_01297_),
    .B2(_01298_),
    .Y(_01299_));
 sky130_fd_sc_hd__or4_1 _05412_ (.A(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .C(_01182_),
    .D(_01195_),
    .X(_01300_));
 sky130_fd_sc_hd__o21a_1 _05413_ (.A1(_01299_),
    .A2(_01300_),
    .B1(_00650_),
    .X(_00648_));
 sky130_fd_sc_hd__nor2_1 _05414_ (.A(_01179_),
    .B(_01196_),
    .Y(_00647_));
 sky130_fd_sc_hd__o21ba_1 _05415_ (.A1(_01236_),
    .A2(net570),
    .B1_N(_01221_),
    .X(_00700_));
 sky130_fd_sc_hd__or3b_1 _05416_ (.A(net731),
    .B(\u_ws281x.u_txd_1.state ),
    .C_N(_01220_),
    .X(_00701_));
 sky130_fd_sc_hd__or2_1 _05417_ (.A(_00826_),
    .B(\u_ws281x.cfg_th1_period[0] ),
    .X(_01301_));
 sky130_fd_sc_hd__and2b_1 _05418_ (.A_N(\u_ws281x.cfg_th1_period[9] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .X(_01302_));
 sky130_fd_sc_hd__a221o_1 _05419_ (.A1(_00826_),
    .A2(\u_ws281x.cfg_th1_period[0] ),
    .B1(_00855_),
    .B2(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .C1(_01302_),
    .X(_01303_));
 sky130_fd_sc_hd__a22o_1 _05420_ (.A1(_00827_),
    .A2(\u_ws281x.cfg_th1_period[1] ),
    .B1(_01301_),
    .B2(_01303_),
    .X(_01304_));
 sky130_fd_sc_hd__o221a_1 _05421_ (.A1(_00827_),
    .A2(\u_ws281x.cfg_th1_period[1] ),
    .B1(\u_ws281x.cfg_th1_period[2] ),
    .B2(_00828_),
    .C1(_01304_),
    .X(_01305_));
 sky130_fd_sc_hd__a21oi_1 _05422_ (.A1(_00828_),
    .A2(\u_ws281x.cfg_th1_period[2] ),
    .B1(_01305_),
    .Y(_01306_));
 sky130_fd_sc_hd__a21oi_1 _05423_ (.A1(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .A2(_00854_),
    .B1(_01306_),
    .Y(_01307_));
 sky130_fd_sc_hd__a22o_1 _05424_ (.A1(_00829_),
    .A2(\u_ws281x.cfg_th1_period[3] ),
    .B1(\u_ws281x.cfg_th1_period[4] ),
    .B2(_00830_),
    .X(_01308_));
 sky130_fd_sc_hd__o22a_1 _05425_ (.A1(_00830_),
    .A2(\u_ws281x.cfg_th1_period[4] ),
    .B1(_01307_),
    .B2(_01308_),
    .X(_01309_));
 sky130_fd_sc_hd__a21o_1 _05426_ (.A1(_00831_),
    .A2(\u_ws281x.cfg_th1_period[5] ),
    .B1(_01309_),
    .X(_01310_));
 sky130_fd_sc_hd__o221a_1 _05427_ (.A1(_00832_),
    .A2(\u_ws281x.cfg_th1_period[6] ),
    .B1(\u_ws281x.cfg_th1_period[5] ),
    .B2(_00831_),
    .C1(_01310_),
    .X(_01311_));
 sky130_fd_sc_hd__a221o_1 _05428_ (.A1(_00833_),
    .A2(\u_ws281x.cfg_th1_period[7] ),
    .B1(\u_ws281x.cfg_th1_period[6] ),
    .B2(_00832_),
    .C1(_01311_),
    .X(_01312_));
 sky130_fd_sc_hd__o221a_1 _05429_ (.A1(_00833_),
    .A2(\u_ws281x.cfg_th1_period[7] ),
    .B1(\u_ws281x.cfg_th1_period[8] ),
    .B2(_00834_),
    .C1(_01312_),
    .X(_01313_));
 sky130_fd_sc_hd__a22o_1 _05430_ (.A1(_00835_),
    .A2(\u_ws281x.cfg_th1_period[9] ),
    .B1(\u_ws281x.cfg_th1_period[8] ),
    .B2(_00834_),
    .X(_01314_));
 sky130_fd_sc_hd__o221a_1 _05431_ (.A1(_00835_),
    .A2(\u_ws281x.cfg_th1_period[9] ),
    .B1(_01313_),
    .B2(_01314_),
    .C1(\u_ws281x.u_txd_1.led_data[23] ),
    .X(_01315_));
 sky130_fd_sc_hd__o211a_1 _05432_ (.A1(_00826_),
    .A2(\u_ws281x.cfg_th0_period[0] ),
    .B1(_00853_),
    .C1(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .X(_01316_));
 sky130_fd_sc_hd__a221o_1 _05433_ (.A1(_00827_),
    .A2(\u_ws281x.cfg_th0_period[1] ),
    .B1(\u_ws281x.cfg_th0_period[0] ),
    .B2(_00826_),
    .C1(_01316_),
    .X(_01317_));
 sky130_fd_sc_hd__o221a_1 _05434_ (.A1(_00828_),
    .A2(\u_ws281x.cfg_th0_period[2] ),
    .B1(\u_ws281x.cfg_th0_period[1] ),
    .B2(_00827_),
    .C1(_01317_),
    .X(_01318_));
 sky130_fd_sc_hd__a221o_1 _05435_ (.A1(_00829_),
    .A2(\u_ws281x.cfg_th0_period[3] ),
    .B1(\u_ws281x.cfg_th0_period[2] ),
    .B2(_00828_),
    .C1(_01318_),
    .X(_01319_));
 sky130_fd_sc_hd__o221a_1 _05436_ (.A1(_00830_),
    .A2(\u_ws281x.cfg_th0_period[4] ),
    .B1(\u_ws281x.cfg_th0_period[3] ),
    .B2(_00829_),
    .C1(_01319_),
    .X(_01320_));
 sky130_fd_sc_hd__a221o_1 _05437_ (.A1(_00831_),
    .A2(\u_ws281x.cfg_th0_period[5] ),
    .B1(\u_ws281x.cfg_th0_period[4] ),
    .B2(_00830_),
    .C1(_01320_),
    .X(_01321_));
 sky130_fd_sc_hd__o221a_1 _05438_ (.A1(_00832_),
    .A2(\u_ws281x.cfg_th0_period[6] ),
    .B1(\u_ws281x.cfg_th0_period[5] ),
    .B2(_00831_),
    .C1(_01321_),
    .X(_01322_));
 sky130_fd_sc_hd__a221o_1 _05439_ (.A1(_00833_),
    .A2(\u_ws281x.cfg_th0_period[7] ),
    .B1(\u_ws281x.cfg_th0_period[6] ),
    .B2(_00832_),
    .C1(_01322_),
    .X(_01323_));
 sky130_fd_sc_hd__o221a_1 _05440_ (.A1(_00834_),
    .A2(\u_ws281x.cfg_th0_period[8] ),
    .B1(\u_ws281x.cfg_th0_period[7] ),
    .B2(_00833_),
    .C1(_01323_),
    .X(_01324_));
 sky130_fd_sc_hd__a221o_1 _05441_ (.A1(_00835_),
    .A2(\u_ws281x.cfg_th0_period[9] ),
    .B1(\u_ws281x.cfg_th0_period[8] ),
    .B2(_00834_),
    .C1(_01324_),
    .X(_01325_));
 sky130_fd_sc_hd__a21oi_1 _05442_ (.A1(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .A2(_00853_),
    .B1(\u_ws281x.u_txd_1.led_data[23] ),
    .Y(_01326_));
 sky130_fd_sc_hd__a21oi_1 _05443_ (.A1(_01325_),
    .A2(_01326_),
    .B1(_01315_),
    .Y(_01327_));
 sky130_fd_sc_hd__or4_1 _05444_ (.A(\u_ws281x.u_txd_1.clk_cnt[11] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[10] ),
    .C(_01223_),
    .D(_01237_),
    .X(_01328_));
 sky130_fd_sc_hd__o21a_1 _05445_ (.A1(_01327_),
    .A2(_01328_),
    .B1(_00701_),
    .X(_00699_));
 sky130_fd_sc_hd__a21oi_1 _05446_ (.A1(\u_ws281x.u_txd_1.state ),
    .A2(_01236_),
    .B1(_01221_),
    .Y(_00698_));
 sky130_fd_sc_hd__or3_1 _05447_ (.A(\u_timer.u_pulse_1ms.cnt[6] ),
    .B(\u_timer.u_pulse_1ms.cnt[9] ),
    .C(\u_timer.u_pulse_1ms.cnt[8] ),
    .X(_01329_));
 sky130_fd_sc_hd__or4_1 _05448_ (.A(\u_timer.u_pulse_1ms.cnt[3] ),
    .B(\u_timer.u_pulse_1ms.cnt[5] ),
    .C(\u_timer.u_pulse_1ms.cnt[4] ),
    .D(\u_timer.u_pulse_1ms.cnt[7] ),
    .X(_01330_));
 sky130_fd_sc_hd__or4b_1 _05449_ (.A(\u_timer.u_pulse_1ms.cnt[1] ),
    .B(\u_timer.u_pulse_1ms.cnt[0] ),
    .C(\u_timer.u_pulse_1ms.cnt[2] ),
    .D_N(\u_gpio.pulse_1us ),
    .X(_01331_));
 sky130_fd_sc_hd__or3_4 _05450_ (.A(_01329_),
    .B(_01330_),
    .C(_01331_),
    .X(_01332_));
 sky130_fd_sc_hd__inv_2 _05451_ (.A(_01332_),
    .Y(net366));
 sky130_fd_sc_hd__and3_1 _05452_ (.A(net1307),
    .B(net1342),
    .C(_01003_),
    .X(_01333_));
 sky130_fd_sc_hd__and3_1 _05453_ (.A(net1416),
    .B(net1341),
    .C(_01333_),
    .X(_01334_));
 sky130_fd_sc_hd__nand3_1 _05454_ (.A(\u_timer.reg_ack ),
    .B(net1180),
    .C(net678),
    .Y(_01335_));
 sky130_fd_sc_hd__nor2_1 _05455_ (.A(\u_timer.cfg_timer0[18] ),
    .B(\u_timer.cfg_timer0[17] ),
    .Y(_01336_));
 sky130_fd_sc_hd__or4_1 _05456_ (.A(\u_timer.u_pulse_1s.cnt[7] ),
    .B(\u_timer.u_pulse_1s.cnt[6] ),
    .C(\u_timer.u_pulse_1s.cnt[9] ),
    .D(\u_timer.u_pulse_1s.cnt[8] ),
    .X(_01337_));
 sky130_fd_sc_hd__or2_1 _05457_ (.A(\u_timer.u_pulse_1s.cnt[1] ),
    .B(\u_timer.u_pulse_1s.cnt[0] ),
    .X(_01338_));
 sky130_fd_sc_hd__or4_1 _05458_ (.A(\u_timer.u_pulse_1s.cnt[3] ),
    .B(\u_timer.u_pulse_1s.cnt[2] ),
    .C(\u_timer.u_pulse_1s.cnt[5] ),
    .D(\u_timer.u_pulse_1s.cnt[4] ),
    .X(_01339_));
 sky130_fd_sc_hd__or3_1 _05459_ (.A(_01337_),
    .B(_01338_),
    .C(_01339_),
    .X(_01340_));
 sky130_fd_sc_hd__a211oi_1 _05460_ (.A1(\u_timer.cfg_timer0[18] ),
    .A2(net567),
    .B1(_01336_),
    .C1(_01332_),
    .Y(_01341_));
 sky130_fd_sc_hd__a21oi_1 _05461_ (.A1(\u_gpio.pulse_1us ),
    .A2(_01336_),
    .B1(_01341_),
    .Y(_01342_));
 sky130_fd_sc_hd__o31a_1 _05462_ (.A1(\u_timer.u_timer_0.timer_counter[15] ),
    .A2(_01268_),
    .A3(_01342_),
    .B1(_01335_),
    .X(_01343_));
 sky130_fd_sc_hd__o21ai_1 _05463_ (.A1(_00848_),
    .A2(_01342_),
    .B1(net521),
    .Y(_00543_));
 sky130_fd_sc_hd__nand3_1 _05464_ (.A(\u_timer.reg_ack ),
    .B(net1160),
    .C(net678),
    .Y(_01344_));
 sky130_fd_sc_hd__or2_1 _05465_ (.A(\u_timer.cfg_timer1[18] ),
    .B(\u_timer.cfg_timer1[17] ),
    .X(_01345_));
 sky130_fd_sc_hd__a2bb2o_1 _05466_ (.A1_N(\u_gpio.pulse_1us ),
    .A2_N(_01345_),
    .B1(net567),
    .B2(\u_timer.cfg_timer1[18] ),
    .X(_01346_));
 sky130_fd_sc_hd__a21o_1 _05467_ (.A1(_01332_),
    .A2(_01345_),
    .B1(_01346_),
    .X(_01347_));
 sky130_fd_sc_hd__o31a_1 _05468_ (.A1(\u_timer.u_timer_1.timer_counter[15] ),
    .A2(_01259_),
    .A3(_01347_),
    .B1(_01344_),
    .X(_01348_));
 sky130_fd_sc_hd__o21ai_1 _05469_ (.A1(_00845_),
    .A2(_01347_),
    .B1(net519),
    .Y(_00560_));
 sky130_fd_sc_hd__nor2_4 _05470_ (.A(net1269),
    .B(net1256),
    .Y(_01349_));
 sky130_fd_sc_hd__nand2_1 _05471_ (.A(net1349),
    .B(net1362),
    .Y(_01350_));
 sky130_fd_sc_hd__or2_1 _05472_ (.A(\u_timer.cfg_timer2[18] ),
    .B(\u_timer.cfg_timer2[17] ),
    .X(_01351_));
 sky130_fd_sc_hd__a2bb2o_1 _05473_ (.A1_N(\u_gpio.pulse_1us ),
    .A2_N(_01351_),
    .B1(net567),
    .B2(\u_timer.cfg_timer2[18] ),
    .X(_01352_));
 sky130_fd_sc_hd__a21o_1 _05474_ (.A1(_01332_),
    .A2(_01351_),
    .B1(_01352_),
    .X(_01353_));
 sky130_fd_sc_hd__nor3_1 _05475_ (.A(\u_timer.u_timer_2.timer_counter[15] ),
    .B(_01250_),
    .C(_01353_),
    .Y(_01354_));
 sky130_fd_sc_hd__a31oi_2 _05476_ (.A1(\u_timer.reg_ack ),
    .A2(net678),
    .A3(net1150),
    .B1(_01354_),
    .Y(_01355_));
 sky130_fd_sc_hd__o21ai_1 _05477_ (.A1(_00842_),
    .A2(_01353_),
    .B1(net515),
    .Y(_00577_));
 sky130_fd_sc_hd__and3_1 _05478_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .C(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .X(_01356_));
 sky130_fd_sc_hd__and2_1 _05479_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ),
    .B(_01356_),
    .X(_01357_));
 sky130_fd_sc_hd__and3_1 _05480_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .C(_01357_),
    .X(_01358_));
 sky130_fd_sc_hd__and2_1 _05481_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ),
    .B(_01358_),
    .X(_01359_));
 sky130_fd_sc_hd__and2_1 _05482_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .B(_01359_),
    .X(_01360_));
 sky130_fd_sc_hd__and3_1 _05483_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .C(_01359_),
    .X(_01361_));
 sky130_fd_sc_hd__and2_1 _05484_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .B(_01361_),
    .X(_01362_));
 sky130_fd_sc_hd__and3_1 _05485_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .C(_01362_),
    .X(_01363_));
 sky130_fd_sc_hd__and2_1 _05486_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .B(_01363_),
    .X(_01364_));
 sky130_fd_sc_hd__and3_1 _05487_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .C(_01364_),
    .X(_01365_));
 sky130_fd_sc_hd__a2bb2o_1 _05488_ (.A1_N(_00866_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_period[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[1] ),
    .B2(_00872_),
    .X(_01366_));
 sky130_fd_sc_hd__a22o_1 _05489_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[5] ),
    .B1(_00876_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .X(_01367_));
 sky130_fd_sc_hd__a221o_1 _05490_ (.A1(_00873_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[0] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[8] ),
    .B2(_00865_),
    .C1(_01367_),
    .X(_01368_));
 sky130_fd_sc_hd__a2bb2o_1 _05491_ (.A1_N(_00865_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_period[8] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[2] ),
    .B2(_00871_),
    .X(_01369_));
 sky130_fd_sc_hd__a221o_1 _05492_ (.A1(net728),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[6] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[7] ),
    .B2(_00866_),
    .C1(_01369_),
    .X(_01370_));
 sky130_fd_sc_hd__a211o_1 _05493_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .A2(_00877_),
    .B1(_01368_),
    .C1(_01370_),
    .X(_01371_));
 sky130_fd_sc_hd__a221o_1 _05494_ (.A1(_00870_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[3] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[15] ),
    .B2(_00858_),
    .C1(_01371_),
    .X(_01372_));
 sky130_fd_sc_hd__o22a_1 _05495_ (.A1(_00863_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[10] ),
    .B1(_00876_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .X(_01373_));
 sky130_fd_sc_hd__xnor2_1 _05496_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_period[9] ),
    .Y(_01374_));
 sky130_fd_sc_hd__a2bb2o_1 _05497_ (.A1_N(_00871_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_period[2] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[4] ),
    .B2(_00869_),
    .X(_01375_));
 sky130_fd_sc_hd__o22ai_1 _05498_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[5] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[6] ),
    .B2(net728),
    .Y(_01376_));
 sky130_fd_sc_hd__o221a_1 _05499_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[4] ),
    .B2(_00869_),
    .C1(_01373_),
    .X(_01377_));
 sky130_fd_sc_hd__o211a_1 _05500_ (.A1(_00873_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[0] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_zeropd ),
    .C1(_01377_),
    .X(_01378_));
 sky130_fd_sc_hd__a221o_1 _05501_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ),
    .A2(_00874_),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[10] ),
    .B2(_00863_),
    .C1(_01376_),
    .X(_01379_));
 sky130_fd_sc_hd__o221ai_1 _05502_ (.A1(_00859_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[14] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[15] ),
    .B2(_00858_),
    .C1(_01374_),
    .Y(_01380_));
 sky130_fd_sc_hd__a221o_1 _05503_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .A2(_00875_),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[14] ),
    .B2(_00859_),
    .C1(_01366_),
    .X(_01381_));
 sky130_fd_sc_hd__a221o_1 _05504_ (.A1(_00862_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_period[11] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_period[13] ),
    .B2(_00860_),
    .C1(_01375_),
    .X(_01382_));
 sky130_fd_sc_hd__or4_1 _05505_ (.A(_01379_),
    .B(_01380_),
    .C(_01381_),
    .D(_01382_),
    .X(_01383_));
 sky130_fd_sc_hd__nor2_1 _05506_ (.A(_01372_),
    .B(_01383_),
    .Y(_01384_));
 sky130_fd_sc_hd__a22o_1 _05507_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[15] ),
    .A2(_01365_),
    .B1(_01378_),
    .B2(_01384_),
    .X(_01385_));
 sky130_fd_sc_hd__nand2_2 _05508_ (.A(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .B(_01385_),
    .Y(_01386_));
 sky130_fd_sc_hd__inv_2 _05509_ (.A(_01386_),
    .Y(\u_pwm.u_pwm_0.u_pwm.pwm_ovflow ));
 sky130_fd_sc_hd__nor2_2 _05510_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_ovflow_l ),
    .B(_01386_),
    .Y(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__inv_2 _05511_ (.A(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .Y(_01387_));
 sky130_fd_sc_hd__nand4b_4 _05512_ (.A_N(net1342),
    .B(_01003_),
    .C(net1307),
    .D(net1341),
    .Y(_01388_));
 sky130_fd_sc_hd__inv_2 _05513_ (.A(_01388_),
    .Y(_01389_));
 sky130_fd_sc_hd__and4_1 _05514_ (.A(net130),
    .B(net1255),
    .C(net1214),
    .D(_01389_),
    .X(_01390_));
 sky130_fd_sc_hd__and4_1 _05515_ (.A(net1334),
    .B(\u_pwm.reg_ack_glbl ),
    .C(net1151),
    .D(_01390_),
    .X(_01391_));
 sky130_fd_sc_hd__a21o_1 _05516_ (.A1(net1296),
    .A2(_01391_),
    .B1(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .X(_00314_));
 sky130_fd_sc_hd__nand2_1 _05517_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .Y(_01392_));
 sky130_fd_sc_hd__nor2_1 _05518_ (.A(_00891_),
    .B(_01392_),
    .Y(_01393_));
 sky130_fd_sc_hd__and4_1 _05519_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .C(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .D(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .X(_01394_));
 sky130_fd_sc_hd__nand2_1 _05520_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .B(_01394_),
    .Y(_01395_));
 sky130_fd_sc_hd__and3_1 _05521_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[5] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .C(_01394_),
    .X(_01396_));
 sky130_fd_sc_hd__and2_1 _05522_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ),
    .B(_01396_),
    .X(_01397_));
 sky130_fd_sc_hd__nand2_1 _05523_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ),
    .B(_01397_),
    .Y(_01398_));
 sky130_fd_sc_hd__and3_1 _05524_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ),
    .C(_01397_),
    .X(_01399_));
 sky130_fd_sc_hd__and2_1 _05525_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .B(_01399_),
    .X(_01400_));
 sky130_fd_sc_hd__nand2_1 _05526_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .B(_01400_),
    .Y(_01401_));
 sky130_fd_sc_hd__and3_1 _05527_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .C(_01400_),
    .X(_01402_));
 sky130_fd_sc_hd__and2_1 _05528_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .B(_01402_),
    .X(_01403_));
 sky130_fd_sc_hd__nand2_1 _05529_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .B(_01403_),
    .Y(_01404_));
 sky130_fd_sc_hd__and3_1 _05530_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .C(_01403_),
    .X(_01405_));
 sky130_fd_sc_hd__o2bb2a_1 _05531_ (.A1_N(_00889_),
    .A2_N(\u_pwm.u_pwm_1.cfg_pwm_period[4] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[12] ),
    .B2(_00881_),
    .X(_01406_));
 sky130_fd_sc_hd__a22oi_1 _05532_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[6] ),
    .B2(_00887_),
    .Y(_01407_));
 sky130_fd_sc_hd__o221a_1 _05533_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .A2(_00894_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[6] ),
    .B2(_00887_),
    .C1(_01407_),
    .X(_01408_));
 sky130_fd_sc_hd__xnor2_1 _05534_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_period[2] ),
    .Y(_01409_));
 sky130_fd_sc_hd__o221a_1 _05535_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .A2(_00896_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[4] ),
    .B2(_00889_),
    .C1(_01409_),
    .X(_01410_));
 sky130_fd_sc_hd__o2111a_1 _05536_ (.A1(_00890_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[3] ),
    .B1(_01406_),
    .C1(_01408_),
    .D1(_01410_),
    .X(_01411_));
 sky130_fd_sc_hd__xnor2_1 _05537_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_period[13] ),
    .Y(_01412_));
 sky130_fd_sc_hd__nor2_1 _05538_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_period[9] ),
    .Y(_01413_));
 sky130_fd_sc_hd__and2_1 _05539_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_period[9] ),
    .X(_01414_));
 sky130_fd_sc_hd__o221a_1 _05540_ (.A1(_00882_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[11] ),
    .B1(_01413_),
    .B2(_01414_),
    .C1(\u_pwm.u_pwm_1.cfg_pwm_zeropd ),
    .X(_01415_));
 sky130_fd_sc_hd__a22o_1 _05541_ (.A1(_00883_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[10] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[15] ),
    .B2(_00878_),
    .X(_01416_));
 sky130_fd_sc_hd__a221o_1 _05542_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .A2(_00894_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[14] ),
    .B2(_00879_),
    .C1(_01416_),
    .X(_01417_));
 sky130_fd_sc_hd__o2bb2a_1 _05543_ (.A1_N(_00881_),
    .A2_N(\u_pwm.u_pwm_1.cfg_pwm_period[12] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[7] ),
    .B2(_00886_),
    .X(_01418_));
 sky130_fd_sc_hd__o221a_1 _05544_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[14] ),
    .B2(_00879_),
    .C1(_01418_),
    .X(_01419_));
 sky130_fd_sc_hd__a22oi_1 _05545_ (.A1(_00886_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[7] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[8] ),
    .B2(_00885_),
    .Y(_01420_));
 sky130_fd_sc_hd__o221a_1 _05546_ (.A1(_00892_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[1] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[8] ),
    .B2(_00885_),
    .C1(_01420_),
    .X(_01421_));
 sky130_fd_sc_hd__o22a_1 _05547_ (.A1(_00883_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_period[10] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_period[15] ),
    .B2(net727),
    .X(_01422_));
 sky130_fd_sc_hd__o221a_1 _05548_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .A2(_00895_),
    .B1(_00897_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .C1(_01422_),
    .X(_01423_));
 sky130_fd_sc_hd__and4b_1 _05549_ (.A_N(_01417_),
    .B(_01419_),
    .C(_01421_),
    .D(_01423_),
    .X(_01424_));
 sky130_fd_sc_hd__and3_1 _05550_ (.A(_01412_),
    .B(_01415_),
    .C(_01424_),
    .X(_01425_));
 sky130_fd_sc_hd__a22o_1 _05551_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ),
    .A2(_01405_),
    .B1(_01411_),
    .B2(_01425_),
    .X(_01426_));
 sky130_fd_sc_hd__nand2_1 _05552_ (.A(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .B(_01426_),
    .Y(_01427_));
 sky130_fd_sc_hd__inv_2 _05553_ (.A(_01427_),
    .Y(\u_pwm.u_pwm_1.u_pwm.pwm_ovflow ));
 sky130_fd_sc_hd__nor2_2 _05554_ (.A(net2190),
    .B(_01427_),
    .Y(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__inv_2 _05555_ (.A(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .Y(_01428_));
 sky130_fd_sc_hd__a21o_1 _05556_ (.A1(net1574),
    .A2(_01391_),
    .B1(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .X(_00315_));
 sky130_fd_sc_hd__nand2_1 _05557_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ),
    .Y(_01429_));
 sky130_fd_sc_hd__nor2_1 _05558_ (.A(net725),
    .B(_01429_),
    .Y(_01430_));
 sky130_fd_sc_hd__and4_1 _05559_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ),
    .C(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .D(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ),
    .X(_01431_));
 sky130_fd_sc_hd__and3_1 _05560_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .C(_01431_),
    .X(_01432_));
 sky130_fd_sc_hd__and2_1 _05561_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .B(_01432_),
    .X(_01433_));
 sky130_fd_sc_hd__and3_1 _05562_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .C(_01432_),
    .X(_01434_));
 sky130_fd_sc_hd__and3_1 _05563_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .C(_01433_),
    .X(_01435_));
 sky130_fd_sc_hd__and2_1 _05564_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .B(_01435_),
    .X(_01436_));
 sky130_fd_sc_hd__and3_1 _05565_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .B(net1073),
    .C(_01436_),
    .X(_01437_));
 sky130_fd_sc_hd__and2_1 _05566_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .B(_01437_),
    .X(_01438_));
 sky130_fd_sc_hd__and3_1 _05567_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .C(_01437_),
    .X(_01439_));
 sky130_fd_sc_hd__or2_1 _05568_ (.A(_00899_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_period[14] ),
    .X(_01440_));
 sky130_fd_sc_hd__xnor2_1 _05569_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_period[9] ),
    .Y(_01441_));
 sky130_fd_sc_hd__o22a_1 _05570_ (.A1(_00913_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[0] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[4] ),
    .B2(_00909_),
    .X(_01442_));
 sky130_fd_sc_hd__o2bb2a_1 _05571_ (.A1_N(_00903_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_period[10] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[15] ),
    .B2(_00898_),
    .X(_01443_));
 sky130_fd_sc_hd__o211ai_1 _05572_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[3] ),
    .B1(_01442_),
    .C1(_01443_),
    .Y(_01444_));
 sky130_fd_sc_hd__a2bb2o_1 _05573_ (.A1_N(_00906_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_period[7] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[1] ),
    .B2(_00912_),
    .X(_01445_));
 sky130_fd_sc_hd__a22o_1 _05574_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .A2(_00915_),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[13] ),
    .B2(_00900_),
    .X(_01446_));
 sky130_fd_sc_hd__a211o_1 _05575_ (.A1(_00899_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[14] ),
    .B1(_01445_),
    .C1(_01446_),
    .X(_01447_));
 sky130_fd_sc_hd__a22o_1 _05576_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[5] ),
    .B1(_00916_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .X(_01448_));
 sky130_fd_sc_hd__a221o_1 _05577_ (.A1(_00913_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[0] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[8] ),
    .B2(_00905_),
    .C1(_01448_),
    .X(_01449_));
 sky130_fd_sc_hd__a2bb2o_1 _05578_ (.A1_N(_00905_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_period[8] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[2] ),
    .B2(_00911_),
    .X(_01450_));
 sky130_fd_sc_hd__a221o_1 _05579_ (.A1(_00907_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[6] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[7] ),
    .B2(_00906_),
    .C1(_01450_),
    .X(_01451_));
 sky130_fd_sc_hd__a211o_1 _05580_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .A2(_00917_),
    .B1(_01449_),
    .C1(_01451_),
    .X(_01452_));
 sky130_fd_sc_hd__a221o_1 _05581_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[3] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[15] ),
    .B2(_00898_),
    .C1(_01452_),
    .X(_01453_));
 sky130_fd_sc_hd__o221a_1 _05582_ (.A1(_00903_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[10] ),
    .B1(_00916_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .C1(_01441_),
    .X(_01454_));
 sky130_fd_sc_hd__o211a_1 _05583_ (.A1(_00912_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[1] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_zeropd ),
    .C1(_01454_),
    .X(_01455_));
 sky130_fd_sc_hd__o22a_1 _05584_ (.A1(net725),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[2] ),
    .B1(_00914_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .X(_01456_));
 sky130_fd_sc_hd__o221a_1 _05585_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_period[5] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_period[6] ),
    .B2(_00907_),
    .C1(_01440_),
    .X(_01457_));
 sky130_fd_sc_hd__o2111a_1 _05586_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .A2(_00915_),
    .B1(_01455_),
    .C1(_01456_),
    .D1(_01457_),
    .X(_01458_));
 sky130_fd_sc_hd__nor4b_1 _05587_ (.A(_01444_),
    .B(_01447_),
    .C(_01453_),
    .D_N(_01458_),
    .Y(_01459_));
 sky130_fd_sc_hd__a31o_1 _05588_ (.A1(net1070),
    .A2(net1072),
    .A3(_01439_),
    .B1(_01459_),
    .X(_01460_));
 sky130_fd_sc_hd__nand2_1 _05589_ (.A(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .B(_01460_),
    .Y(_01461_));
 sky130_fd_sc_hd__clkinv_2 _05590_ (.A(_01461_),
    .Y(\u_pwm.u_pwm_2.u_pwm.pwm_ovflow ));
 sky130_fd_sc_hd__nor2_4 _05591_ (.A(net2341),
    .B(_01461_),
    .Y(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ));
 sky130_fd_sc_hd__inv_2 _05592_ (.A(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .Y(_01462_));
 sky130_fd_sc_hd__a21o_1 _05593_ (.A1(net1490),
    .A2(_01391_),
    .B1(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .X(_00316_));
 sky130_fd_sc_hd__a21oi_1 _05594_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .A2(_01387_),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_dupdate ),
    .Y(_00353_));
 sky130_fd_sc_hd__and3b_1 _05595_ (.A_N(\u_pwm.u_pwm_0.gpio_tgr ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_run ),
    .C(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .X(_01463_));
 sky130_fd_sc_hd__and2_1 _05596_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ),
    .X(_01464_));
 sky130_fd_sc_hd__and3_1 _05597_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[3] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ),
    .C(_01464_),
    .X(_01465_));
 sky130_fd_sc_hd__o21a_1 _05598_ (.A1(_00919_),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[5] ),
    .X(_01466_));
 sky130_fd_sc_hd__nor2_1 _05599_ (.A(\u_pwm.u_pwm_0.cfg_pwm_scale[0] ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_scale[1] ),
    .Y(_01467_));
 sky130_fd_sc_hd__o21ai_1 _05600_ (.A1(_00919_),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ),
    .Y(_01468_));
 sky130_fd_sc_hd__a2bb2o_1 _05601_ (.A1_N(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ),
    .A2_N(_01467_),
    .B1(_01468_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_scale[1] ),
    .X(_01469_));
 sky130_fd_sc_hd__o21ai_1 _05602_ (.A1(_00920_),
    .A2(_01466_),
    .B1(_01465_),
    .Y(_01470_));
 sky130_fd_sc_hd__o21ai_1 _05603_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ),
    .A2(_01467_),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_scale[2] ),
    .Y(_01471_));
 sky130_fd_sc_hd__o22a_1 _05604_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_scale[2] ),
    .A2(_01469_),
    .B1(_01470_),
    .B2(_01471_),
    .X(_01472_));
 sky130_fd_sc_hd__o21ai_1 _05605_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_scale[3] ),
    .A2(_01472_),
    .B1(net676),
    .Y(_01473_));
 sky130_fd_sc_hd__and3_1 _05606_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[5] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ),
    .C(_01465_),
    .X(_01474_));
 sky130_fd_sc_hd__and3_1 _05607_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[7] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ),
    .C(_01474_),
    .X(_01475_));
 sky130_fd_sc_hd__o21a_1 _05608_ (.A1(_00919_),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[14] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[13] ),
    .X(_01476_));
 sky130_fd_sc_hd__o221a_1 _05609_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ),
    .A2(_01467_),
    .B1(_01476_),
    .B2(_00920_),
    .C1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[11] ),
    .X(_01477_));
 sky130_fd_sc_hd__or2_1 _05610_ (.A(_00918_),
    .B(_01477_),
    .X(_01478_));
 sky130_fd_sc_hd__a21o_1 _05611_ (.A1(_00918_),
    .A2(_00919_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ),
    .X(_01479_));
 sky130_fd_sc_hd__a22o_1 _05612_ (.A1(_00918_),
    .A2(_00920_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[9] ),
    .B2(_01479_),
    .X(_01480_));
 sky130_fd_sc_hd__a32o_1 _05613_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ),
    .A2(_01478_),
    .A3(_01480_),
    .B1(_01467_),
    .B2(_00918_),
    .X(_01481_));
 sky130_fd_sc_hd__a31o_1 _05614_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_scale[3] ),
    .A2(_01475_),
    .A3(_01481_),
    .B1(_01473_),
    .X(_00350_));
 sky130_fd_sc_hd__nand2b_1 _05615_ (.A_N(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_hold ),
    .Y(_00351_));
 sky130_fd_sc_hd__a21oi_1 _05616_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .A2(_01428_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_dupdate ),
    .Y(_00406_));
 sky130_fd_sc_hd__and3b_2 _05617_ (.A_N(\u_pwm.u_pwm_1.gpio_tgr ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_run ),
    .C(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .X(_01482_));
 sky130_fd_sc_hd__and2_1 _05618_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ),
    .X(_01483_));
 sky130_fd_sc_hd__and3_1 _05619_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[3] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ),
    .C(_01483_),
    .X(_01484_));
 sky130_fd_sc_hd__o21a_1 _05620_ (.A1(_00922_),
    .A2(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[5] ),
    .X(_01485_));
 sky130_fd_sc_hd__nor2_1 _05621_ (.A(\u_pwm.u_pwm_1.cfg_pwm_scale[0] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_scale[1] ),
    .Y(_01486_));
 sky130_fd_sc_hd__o21ai_1 _05622_ (.A1(_00922_),
    .A2(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ),
    .Y(_01487_));
 sky130_fd_sc_hd__a2bb2o_1 _05623_ (.A1_N(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ),
    .A2_N(_01486_),
    .B1(_01487_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_scale[1] ),
    .X(_01488_));
 sky130_fd_sc_hd__o21ai_1 _05624_ (.A1(_00923_),
    .A2(_01485_),
    .B1(_01484_),
    .Y(_01489_));
 sky130_fd_sc_hd__o21ai_1 _05625_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ),
    .A2(_01486_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_scale[2] ),
    .Y(_01490_));
 sky130_fd_sc_hd__o22a_1 _05626_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_scale[2] ),
    .A2(_01488_),
    .B1(_01489_),
    .B2(_01490_),
    .X(_01491_));
 sky130_fd_sc_hd__o21ai_1 _05627_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_scale[3] ),
    .A2(_01491_),
    .B1(net674),
    .Y(_01492_));
 sky130_fd_sc_hd__o21a_1 _05628_ (.A1(_00922_),
    .A2(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[14] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[13] ),
    .X(_01493_));
 sky130_fd_sc_hd__o221a_1 _05629_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ),
    .A2(_01486_),
    .B1(_01493_),
    .B2(_00923_),
    .C1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[11] ),
    .X(_01494_));
 sky130_fd_sc_hd__or2_1 _05630_ (.A(_00921_),
    .B(_01494_),
    .X(_01495_));
 sky130_fd_sc_hd__a21o_1 _05631_ (.A1(_00921_),
    .A2(_00922_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ),
    .X(_01496_));
 sky130_fd_sc_hd__a22o_1 _05632_ (.A1(_00921_),
    .A2(_00923_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[9] ),
    .B2(_01496_),
    .X(_01497_));
 sky130_fd_sc_hd__a32o_1 _05633_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ),
    .A2(_01495_),
    .A3(_01497_),
    .B1(_01486_),
    .B2(_00921_),
    .X(_01498_));
 sky130_fd_sc_hd__and3_1 _05634_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[5] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ),
    .C(_01484_),
    .X(_01499_));
 sky130_fd_sc_hd__and3_1 _05635_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[7] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ),
    .C(_01499_),
    .X(_01500_));
 sky130_fd_sc_hd__a31o_1 _05636_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_scale[3] ),
    .A2(_01498_),
    .A3(_01500_),
    .B1(_01492_),
    .X(_00403_));
 sky130_fd_sc_hd__nand2b_1 _05637_ (.A_N(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_hold ),
    .Y(_00404_));
 sky130_fd_sc_hd__a21oi_4 _05638_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .A2(_01462_),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_dupdate ),
    .Y(_00459_));
 sky130_fd_sc_hd__and3b_1 _05639_ (.A_N(\u_pwm.u_pwm_2.gpio_tgr ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_run ),
    .C(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .X(_01501_));
 sky130_fd_sc_hd__and2_1 _05640_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ),
    .X(_01502_));
 sky130_fd_sc_hd__and3_1 _05641_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[3] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ),
    .C(_01502_),
    .X(_01503_));
 sky130_fd_sc_hd__o21a_1 _05642_ (.A1(_00925_),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[5] ),
    .X(_01504_));
 sky130_fd_sc_hd__nor2_1 _05643_ (.A(\u_pwm.u_pwm_2.cfg_pwm_scale[0] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_scale[1] ),
    .Y(_01505_));
 sky130_fd_sc_hd__o21ai_1 _05644_ (.A1(_00925_),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ),
    .Y(_01506_));
 sky130_fd_sc_hd__a2bb2o_1 _05645_ (.A1_N(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ),
    .A2_N(_01505_),
    .B1(_01506_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_scale[1] ),
    .X(_01507_));
 sky130_fd_sc_hd__o21ai_1 _05646_ (.A1(_00926_),
    .A2(_01504_),
    .B1(_01503_),
    .Y(_01508_));
 sky130_fd_sc_hd__o21ai_1 _05647_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ),
    .A2(_01505_),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_scale[2] ),
    .Y(_01509_));
 sky130_fd_sc_hd__o22a_1 _05648_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_scale[2] ),
    .A2(_01507_),
    .B1(_01508_),
    .B2(_01509_),
    .X(_01510_));
 sky130_fd_sc_hd__o21ai_1 _05649_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_scale[3] ),
    .A2(_01510_),
    .B1(net672),
    .Y(_01511_));
 sky130_fd_sc_hd__and3_1 _05650_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[5] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ),
    .C(_01503_),
    .X(_01512_));
 sky130_fd_sc_hd__and3_1 _05651_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[7] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ),
    .C(_01512_),
    .X(_01513_));
 sky130_fd_sc_hd__o21a_1 _05652_ (.A1(_00925_),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[14] ),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[13] ),
    .X(_01514_));
 sky130_fd_sc_hd__o221a_1 _05653_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ),
    .A2(_01505_),
    .B1(_01514_),
    .B2(_00926_),
    .C1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[11] ),
    .X(_01515_));
 sky130_fd_sc_hd__or2_1 _05654_ (.A(_00924_),
    .B(_01515_),
    .X(_01516_));
 sky130_fd_sc_hd__a21o_1 _05655_ (.A1(_00924_),
    .A2(_00925_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ),
    .X(_01517_));
 sky130_fd_sc_hd__a22o_1 _05656_ (.A1(_00924_),
    .A2(_00926_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[9] ),
    .B2(_01517_),
    .X(_01518_));
 sky130_fd_sc_hd__a32o_1 _05657_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ),
    .A2(_01516_),
    .A3(_01518_),
    .B1(_01505_),
    .B2(_00924_),
    .X(_01519_));
 sky130_fd_sc_hd__a31o_1 _05658_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_scale[3] ),
    .A2(_01513_),
    .A3(_01519_),
    .B1(_01511_),
    .X(_00456_));
 sky130_fd_sc_hd__nand2b_1 _05659_ (.A_N(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_hold ),
    .Y(_00457_));
 sky130_fd_sc_hd__xor2_1 _05660_ (.A(\u_timer.u_pulse_1us.cnt[5] ),
    .B(\u_timer.cfg_pulse_1us[5] ),
    .X(_01520_));
 sky130_fd_sc_hd__o22ai_1 _05661_ (.A1(\u_timer.u_pulse_1us.cnt[1] ),
    .A2(_00927_),
    .B1(_00928_),
    .B2(\u_timer.cfg_pulse_1us[3] ),
    .Y(_01521_));
 sky130_fd_sc_hd__xnor2_1 _05662_ (.A(\u_timer.u_pulse_1us.cnt[0] ),
    .B(\u_timer.cfg_pulse_1us[0] ),
    .Y(_01522_));
 sky130_fd_sc_hd__o22ai_1 _05663_ (.A1(\u_timer.u_pulse_1us.cnt[4] ),
    .A2(_00929_),
    .B1(_00934_),
    .B2(\u_timer.cfg_pulse_1us[9] ),
    .Y(_01523_));
 sky130_fd_sc_hd__a22o_1 _05664_ (.A1(\u_timer.u_pulse_1us.cnt[1] ),
    .A2(_00927_),
    .B1(_00934_),
    .B2(\u_timer.cfg_pulse_1us[9] ),
    .X(_01524_));
 sky130_fd_sc_hd__xor2_1 _05665_ (.A(\u_timer.u_pulse_1us.cnt[2] ),
    .B(\u_timer.cfg_pulse_1us[2] ),
    .X(_01525_));
 sky130_fd_sc_hd__a22o_1 _05666_ (.A1(_00928_),
    .A2(\u_timer.cfg_pulse_1us[3] ),
    .B1(_00931_),
    .B2(\u_timer.cfg_pulse_1us[7] ),
    .X(_01526_));
 sky130_fd_sc_hd__a221o_1 _05667_ (.A1(\u_timer.u_pulse_1us.cnt[7] ),
    .A2(_00932_),
    .B1(_00933_),
    .B2(\u_timer.cfg_pulse_1us[8] ),
    .C1(_01521_),
    .X(_01527_));
 sky130_fd_sc_hd__o221a_1 _05668_ (.A1(_00930_),
    .A2(\u_timer.cfg_pulse_1us[6] ),
    .B1(_00933_),
    .B2(\u_timer.cfg_pulse_1us[8] ),
    .C1(_01522_),
    .X(_01528_));
 sky130_fd_sc_hd__a221o_1 _05669_ (.A1(\u_timer.u_pulse_1us.cnt[4] ),
    .A2(_00929_),
    .B1(_00930_),
    .B2(\u_timer.cfg_pulse_1us[6] ),
    .C1(_01526_),
    .X(_01529_));
 sky130_fd_sc_hd__or4b_1 _05670_ (.A(_01524_),
    .B(_01529_),
    .C(_01525_),
    .D_N(_01528_),
    .X(_01530_));
 sky130_fd_sc_hd__or4_4 _05671_ (.A(_01520_),
    .B(_01523_),
    .C(_01527_),
    .D(_01530_),
    .X(_01531_));
 sky130_fd_sc_hd__inv_2 _05672_ (.A(_01531_),
    .Y(_00499_));
 sky130_fd_sc_hd__or4_4 _05673_ (.A(_00776_),
    .B(net1344),
    .C(_00997_),
    .D(_01388_),
    .X(_01532_));
 sky130_fd_sc_hd__nor2_2 _05674_ (.A(net1212),
    .B(_01532_),
    .Y(_01533_));
 sky130_fd_sc_hd__and2_1 _05675_ (.A(net1313),
    .B(_01533_),
    .X(_00367_));
 sky130_fd_sc_hd__or4_4 _05676_ (.A(_00776_),
    .B(net1344),
    .C(_01117_),
    .D(_01388_),
    .X(_01534_));
 sky130_fd_sc_hd__nor2_1 _05677_ (.A(net1212),
    .B(_01534_),
    .Y(_01535_));
 sky130_fd_sc_hd__and2_1 _05678_ (.A(net1311),
    .B(_01535_),
    .X(_00420_));
 sky130_fd_sc_hd__or3_4 _05679_ (.A(_00776_),
    .B(_01145_),
    .C(_01388_),
    .X(_01536_));
 sky130_fd_sc_hd__nor2_4 _05680_ (.A(net1211),
    .B(_01536_),
    .Y(_01537_));
 sky130_fd_sc_hd__and2_1 _05681_ (.A(net1310),
    .B(_01537_),
    .X(_00473_));
 sky130_fd_sc_hd__nor2_4 _05682_ (.A(_00997_),
    .B(net1212),
    .Y(_01538_));
 sky130_fd_sc_hd__and3_1 _05683_ (.A(net1310),
    .B(net1175),
    .C(net669),
    .X(_00301_));
 sky130_fd_sc_hd__nor2_2 _05684_ (.A(_00997_),
    .B(_01115_),
    .Y(_01539_));
 sky130_fd_sc_hd__and3_1 _05685_ (.A(net1310),
    .B(net1175),
    .C(net665),
    .X(_00297_));
 sky130_fd_sc_hd__nor2_1 _05686_ (.A(_01130_),
    .B(net1212),
    .Y(_01540_));
 sky130_fd_sc_hd__and3_1 _05687_ (.A(net1310),
    .B(net1175),
    .C(net1136),
    .X(_00261_));
 sky130_fd_sc_hd__and3_1 _05688_ (.A(net1311),
    .B(net1175),
    .C(net702),
    .X(_00257_));
 sky130_fd_sc_hd__nor2_2 _05689_ (.A(net1228),
    .B(_01130_),
    .Y(_01541_));
 sky130_fd_sc_hd__and3_1 _05690_ (.A(net1311),
    .B(net1175),
    .C(net1132),
    .X(_00253_));
 sky130_fd_sc_hd__and4b_1 _05691_ (.A_N(\u_gpio.reg_ack ),
    .B(net1342),
    .C(_01002_),
    .D(_01003_),
    .X(_00251_));
 sky130_fd_sc_hd__nor2_1 _05692_ (.A(net1228),
    .B(_01117_),
    .Y(_01542_));
 sky130_fd_sc_hd__and3_1 _05693_ (.A(net1334),
    .B(net1175),
    .C(net660),
    .X(_00306_));
 sky130_fd_sc_hd__and3_1 _05694_ (.A(net1325),
    .B(net1176),
    .C(net663),
    .X(_00307_));
 sky130_fd_sc_hd__and3_1 _05695_ (.A(net1319),
    .B(net1177),
    .C(net661),
    .X(_00304_));
 sky130_fd_sc_hd__and3_1 _05696_ (.A(net1334),
    .B(net1177),
    .C(net670),
    .X(_00302_));
 sky130_fd_sc_hd__and3_1 _05697_ (.A(net1324),
    .B(net1176),
    .C(net668),
    .X(_00303_));
 sky130_fd_sc_hd__and3_1 _05698_ (.A(net1321),
    .B(net1177),
    .C(net671),
    .X(_00300_));
 sky130_fd_sc_hd__and3_1 _05699_ (.A(net1334),
    .B(net1177),
    .C(net667),
    .X(_00298_));
 sky130_fd_sc_hd__and3_1 _05700_ (.A(net1325),
    .B(net1176),
    .C(net664),
    .X(_00299_));
 sky130_fd_sc_hd__and3_1 _05701_ (.A(net1319),
    .B(net1178),
    .C(net666),
    .X(_00296_));
 sky130_fd_sc_hd__and3_1 _05702_ (.A(net1334),
    .B(net1175),
    .C(net1138),
    .X(_00262_));
 sky130_fd_sc_hd__and3_1 _05703_ (.A(net1325),
    .B(net1176),
    .C(net1137),
    .X(_00263_));
 sky130_fd_sc_hd__and3_1 _05704_ (.A(net1319),
    .B(net1177),
    .C(net1139),
    .X(_00260_));
 sky130_fd_sc_hd__and3_1 _05705_ (.A(net1334),
    .B(net1176),
    .C(net704),
    .X(_00258_));
 sky130_fd_sc_hd__and3_1 _05706_ (.A(net1324),
    .B(net1175),
    .C(net702),
    .X(_00259_));
 sky130_fd_sc_hd__and3_1 _05707_ (.A(net1320),
    .B(net1177),
    .C(net707),
    .X(_00256_));
 sky130_fd_sc_hd__and3_1 _05708_ (.A(net1334),
    .B(net1176),
    .C(net1133),
    .X(_00254_));
 sky130_fd_sc_hd__and3_1 _05709_ (.A(net1324),
    .B(net1175),
    .C(net1131),
    .X(_00255_));
 sky130_fd_sc_hd__and3_1 _05710_ (.A(net1320),
    .B(net1178),
    .C(net1134),
    .X(_00252_));
 sky130_fd_sc_hd__and3_1 _05711_ (.A(net1310),
    .B(net1175),
    .C(net659),
    .X(_00305_));
 sky130_fd_sc_hd__and3_1 _05712_ (.A(net1357),
    .B(net1369),
    .C(_01144_),
    .X(_01543_));
 sky130_fd_sc_hd__nand2_1 _05713_ (.A(_01144_),
    .B(net1145),
    .Y(_01544_));
 sky130_fd_sc_hd__nor2_2 _05714_ (.A(_01145_),
    .B(net1212),
    .Y(_01545_));
 sky130_fd_sc_hd__and3_1 _05715_ (.A(net1319),
    .B(net1173),
    .C(net657),
    .X(_00127_));
 sky130_fd_sc_hd__and3_1 _05716_ (.A(net1324),
    .B(net1169),
    .C(net657),
    .X(_00130_));
 sky130_fd_sc_hd__and3_1 _05717_ (.A(net1331),
    .B(net1167),
    .C(net655),
    .X(_00129_));
 sky130_fd_sc_hd__and3_2 _05718_ (.A(net1343),
    .B(net1247),
    .C(net1214),
    .X(_01546_));
 sky130_fd_sc_hd__and3_1 _05719_ (.A(net1319),
    .B(net1173),
    .C(net1127),
    .X(_00133_));
 sky130_fd_sc_hd__and3_1 _05720_ (.A(net1323),
    .B(net1172),
    .C(net1128),
    .X(_00132_));
 sky130_fd_sc_hd__and3_1 _05721_ (.A(net1332),
    .B(net1168),
    .C(net1124),
    .X(_00131_));
 sky130_fd_sc_hd__and3_1 _05722_ (.A(net1343),
    .B(net1179),
    .C(net1214),
    .X(_01547_));
 sky130_fd_sc_hd__and3_1 _05723_ (.A(net1319),
    .B(net1172),
    .C(net652),
    .X(_00135_));
 sky130_fd_sc_hd__and3_1 _05724_ (.A(net1323),
    .B(net1172),
    .C(net652),
    .X(_00137_));
 sky130_fd_sc_hd__and3_1 _05725_ (.A(net1331),
    .B(net1168),
    .C(net650),
    .X(_00138_));
 sky130_fd_sc_hd__and3_2 _05726_ (.A(net1343),
    .B(net1161),
    .C(net1214),
    .X(_01548_));
 sky130_fd_sc_hd__and3_1 _05727_ (.A(net1316),
    .B(net1169),
    .C(net648),
    .X(_00141_));
 sky130_fd_sc_hd__and3_1 _05728_ (.A(net1323),
    .B(net1172),
    .C(net647),
    .X(_00139_));
 sky130_fd_sc_hd__and3_1 _05729_ (.A(net1331),
    .B(net1167),
    .C(net645),
    .X(_00142_));
 sky130_fd_sc_hd__and2_1 _05730_ (.A(net1343),
    .B(net1139),
    .X(_01549_));
 sky130_fd_sc_hd__and3_1 _05731_ (.A(net1319),
    .B(net1173),
    .C(net644),
    .X(_00143_));
 sky130_fd_sc_hd__and3_1 _05732_ (.A(net1323),
    .B(net1169),
    .C(net643),
    .X(_00146_));
 sky130_fd_sc_hd__and3_1 _05733_ (.A(net1331),
    .B(net1167),
    .C(net641),
    .X(_00145_));
 sky130_fd_sc_hd__and3_4 _05734_ (.A(net1343),
    .B(net1181),
    .C(net1247),
    .X(_01550_));
 sky130_fd_sc_hd__and3_1 _05735_ (.A(net1319),
    .B(net1173),
    .C(net640),
    .X(_00151_));
 sky130_fd_sc_hd__and3_1 _05736_ (.A(net1323),
    .B(net1170),
    .C(net639),
    .X(_00154_));
 sky130_fd_sc_hd__and3_1 _05737_ (.A(net1332),
    .B(net1167),
    .C(net638),
    .X(_00153_));
 sky130_fd_sc_hd__and3_2 _05738_ (.A(net1343),
    .B(net1181),
    .C(net1179),
    .X(_01551_));
 sky130_fd_sc_hd__and3_1 _05739_ (.A(net1319),
    .B(net1172),
    .C(net635),
    .X(_00155_));
 sky130_fd_sc_hd__and3_1 _05740_ (.A(net1323),
    .B(net1172),
    .C(net635),
    .X(_00158_));
 sky130_fd_sc_hd__and3_1 _05741_ (.A(net1332),
    .B(net1168),
    .C(net634),
    .X(_00157_));
 sky130_fd_sc_hd__and3_1 _05742_ (.A(net1343),
    .B(net1181),
    .C(net1160),
    .X(_01552_));
 sky130_fd_sc_hd__and3_1 _05743_ (.A(net1319),
    .B(net1173),
    .C(net631),
    .X(_00159_));
 sky130_fd_sc_hd__and3_1 _05744_ (.A(net1323),
    .B(net1172),
    .C(net630),
    .X(_00162_));
 sky130_fd_sc_hd__and3_1 _05745_ (.A(net1331),
    .B(net1167),
    .C(net629),
    .X(_00161_));
 sky130_fd_sc_hd__and3_4 _05746_ (.A(net1343),
    .B(net1181),
    .C(net1145),
    .X(_01553_));
 sky130_fd_sc_hd__and3_1 _05747_ (.A(net1316),
    .B(net1169),
    .C(net626),
    .X(_00163_));
 sky130_fd_sc_hd__and3_1 _05748_ (.A(net1324),
    .B(net1169),
    .C(net627),
    .X(_00166_));
 sky130_fd_sc_hd__and3_1 _05749_ (.A(net1331),
    .B(net1167),
    .C(net624),
    .X(_00165_));
 sky130_fd_sc_hd__and2_2 _05750_ (.A(net1254),
    .B(net1137),
    .X(_01554_));
 sky130_fd_sc_hd__and3_1 _05751_ (.A(net1316),
    .B(net1173),
    .C(net623),
    .X(_00167_));
 sky130_fd_sc_hd__and3_1 _05752_ (.A(net1324),
    .B(net1170),
    .C(net622),
    .X(_00170_));
 sky130_fd_sc_hd__and3_1 _05753_ (.A(net1335),
    .B(net1170),
    .C(net622),
    .X(_00169_));
 sky130_fd_sc_hd__and3_1 _05754_ (.A(net1254),
    .B(net1181),
    .C(net1179),
    .X(_01555_));
 sky130_fd_sc_hd__and3_1 _05755_ (.A(net1316),
    .B(net1172),
    .C(net618),
    .X(_00173_));
 sky130_fd_sc_hd__and3_1 _05756_ (.A(net1324),
    .B(net1170),
    .C(net617),
    .X(_00172_));
 sky130_fd_sc_hd__and3_1 _05757_ (.A(net1332),
    .B(net1171),
    .C(net617),
    .X(_00171_));
 sky130_fd_sc_hd__and3_1 _05758_ (.A(net1254),
    .B(net1181),
    .C(net1161),
    .X(_01556_));
 sky130_fd_sc_hd__and3_1 _05759_ (.A(net1316),
    .B(net1169),
    .C(net614),
    .X(_00175_));
 sky130_fd_sc_hd__and3_1 _05760_ (.A(net1324),
    .B(net1168),
    .C(net613),
    .X(_00178_));
 sky130_fd_sc_hd__and3_1 _05761_ (.A(net1332),
    .B(net1167),
    .C(net612),
    .X(_00177_));
 sky130_fd_sc_hd__and3_2 _05762_ (.A(net1254),
    .B(net1181),
    .C(net1145),
    .X(_01557_));
 sky130_fd_sc_hd__and3_1 _05763_ (.A(net1317),
    .B(net1169),
    .C(net610),
    .X(_00180_));
 sky130_fd_sc_hd__and3_1 _05764_ (.A(net1323),
    .B(net1169),
    .C(net611),
    .X(_00179_));
 sky130_fd_sc_hd__and3_1 _05765_ (.A(net1331),
    .B(net1167),
    .C(net607),
    .X(_00182_));
 sky130_fd_sc_hd__and3_1 _05766_ (.A(net1255),
    .B(net1247),
    .C(net1153),
    .X(_01558_));
 sky130_fd_sc_hd__and3_1 _05767_ (.A(net1320),
    .B(net1174),
    .C(net605),
    .X(_00185_));
 sky130_fd_sc_hd__and3_1 _05768_ (.A(net1329),
    .B(net1174),
    .C(net606),
    .X(_00184_));
 sky130_fd_sc_hd__and3_1 _05769_ (.A(net1336),
    .B(net1174),
    .C(net606),
    .X(_00183_));
 sky130_fd_sc_hd__and4bb_1 _05770_ (.A_N(net1342),
    .B_N(\u_glbl_reg.reg_ack ),
    .C(_01002_),
    .D(_01003_),
    .X(_00038_));
 sky130_fd_sc_hd__and3_1 _05771_ (.A(net1308),
    .B(net1166),
    .C(net654),
    .X(_00128_));
 sky130_fd_sc_hd__and3_1 _05772_ (.A(net1309),
    .B(net1170),
    .C(net1126),
    .X(_00134_));
 sky130_fd_sc_hd__and3_1 _05773_ (.A(net1309),
    .B(net1168),
    .C(net649),
    .X(_00136_));
 sky130_fd_sc_hd__and3_1 _05774_ (.A(net1308),
    .B(net1166),
    .C(net645),
    .X(_00140_));
 sky130_fd_sc_hd__and3_1 _05775_ (.A(net1309),
    .B(net1168),
    .C(net641),
    .X(_00144_));
 sky130_fd_sc_hd__and3_1 _05776_ (.A(net1308),
    .B(net1166),
    .C(net637),
    .X(_00152_));
 sky130_fd_sc_hd__and3_1 _05777_ (.A(net1308),
    .B(net1166),
    .C(net633),
    .X(_00156_));
 sky130_fd_sc_hd__and3_1 _05778_ (.A(net1309),
    .B(net1168),
    .C(net628),
    .X(_00160_));
 sky130_fd_sc_hd__and3_1 _05779_ (.A(net1308),
    .B(net1166),
    .C(net624),
    .X(_00164_));
 sky130_fd_sc_hd__and3_1 _05780_ (.A(net1309),
    .B(net1168),
    .C(net620),
    .X(_00168_));
 sky130_fd_sc_hd__and3_1 _05781_ (.A(net1308),
    .B(net1166),
    .C(net616),
    .X(_00174_));
 sky130_fd_sc_hd__and3_1 _05782_ (.A(net1309),
    .B(net1168),
    .C(net615),
    .X(_00176_));
 sky130_fd_sc_hd__and3_1 _05783_ (.A(net1309),
    .B(net1168),
    .C(net607),
    .X(_00181_));
 sky130_fd_sc_hd__and3_1 _05784_ (.A(net1313),
    .B(net1174),
    .C(net605),
    .X(_00186_));
 sky130_fd_sc_hd__and2_2 _05785_ (.A(net1216),
    .B(_01270_),
    .X(_01559_));
 sky130_fd_sc_hd__and3_1 _05786_ (.A(net1329),
    .B(net1180),
    .C(_01559_),
    .X(_00594_));
 sky130_fd_sc_hd__nand3b_1 _05787_ (.A_N(\u_ws281x.reg_ack ),
    .B(_01002_),
    .C(_01269_),
    .Y(_01560_));
 sky130_fd_sc_hd__nor2_1 _05788_ (.A(net1416),
    .B(_01560_),
    .Y(_00579_));
 sky130_fd_sc_hd__and3_1 _05789_ (.A(net1337),
    .B(net696),
    .C(_01270_),
    .X(_00598_));
 sky130_fd_sc_hd__and3_1 _05790_ (.A(net1329),
    .B(net1164),
    .C(_01559_),
    .X(_00599_));
 sky130_fd_sc_hd__and3_1 _05791_ (.A(net1322),
    .B(net1165),
    .C(_01559_),
    .X(_00596_));
 sky130_fd_sc_hd__and3_1 _05792_ (.A(net1337),
    .B(net1180),
    .C(_01559_),
    .X(_00595_));
 sky130_fd_sc_hd__and3_1 _05793_ (.A(net1313),
    .B(net1164),
    .C(_01559_),
    .X(_00597_));
 sky130_fd_sc_hd__and3_1 _05794_ (.A(net1311),
    .B(net1159),
    .C(net680),
    .X(_00520_));
 sky130_fd_sc_hd__and3_1 _05795_ (.A(net1314),
    .B(net1179),
    .C(net680),
    .X(_00516_));
 sky130_fd_sc_hd__and3_1 _05796_ (.A(net1311),
    .B(net1247),
    .C(net680),
    .X(_00512_));
 sky130_fd_sc_hd__and3b_1 _05797_ (.A_N(\u_timer.reg_ack ),
    .B(_01333_),
    .C(net1341),
    .X(_00510_));
 sky130_fd_sc_hd__and3_1 _05798_ (.A(net1337),
    .B(net678),
    .C(net1149),
    .X(_00525_));
 sky130_fd_sc_hd__and3_1 _05799_ (.A(net1329),
    .B(net679),
    .C(net1148),
    .X(_00526_));
 sky130_fd_sc_hd__and3_1 _05800_ (.A(net1320),
    .B(net678),
    .C(net1150),
    .X(_00523_));
 sky130_fd_sc_hd__and3_1 _05801_ (.A(net1337),
    .B(net1165),
    .C(net678),
    .X(_00521_));
 sky130_fd_sc_hd__and3_1 _05802_ (.A(net1329),
    .B(net1165),
    .C(net678),
    .X(_00522_));
 sky130_fd_sc_hd__and3_1 _05803_ (.A(net1320),
    .B(net1160),
    .C(net678),
    .X(_00519_));
 sky130_fd_sc_hd__and3_1 _05804_ (.A(net1337),
    .B(net1180),
    .C(net679),
    .X(_00517_));
 sky130_fd_sc_hd__and3_1 _05805_ (.A(net1329),
    .B(net1180),
    .C(net679),
    .X(_00518_));
 sky130_fd_sc_hd__and3_1 _05806_ (.A(net1322),
    .B(net1180),
    .C(net678),
    .X(_00515_));
 sky130_fd_sc_hd__and3_1 _05807_ (.A(net1337),
    .B(net1250),
    .C(net679),
    .X(_00513_));
 sky130_fd_sc_hd__and3_1 _05808_ (.A(net1329),
    .B(net1250),
    .C(net679),
    .X(_00514_));
 sky130_fd_sc_hd__and3_1 _05809_ (.A(net1322),
    .B(net1248),
    .C(net678),
    .X(_00511_));
 sky130_fd_sc_hd__and3_1 _05810_ (.A(net1314),
    .B(net680),
    .C(net1145),
    .X(_00524_));
 sky130_fd_sc_hd__or4bb_1 _05811_ (.A(net1342),
    .B(net1374),
    .C_N(net1340),
    .D_N(_01002_),
    .X(_01561_));
 sky130_fd_sc_hd__o21ai_1 _05812_ (.A1(_00776_),
    .A2(_01561_),
    .B1(net1129),
    .Y(_01562_));
 sky130_fd_sc_hd__o211a_1 _05813_ (.A1(net1336),
    .A2(_01544_),
    .B1(_01562_),
    .C1(\u_semaphore.reg_ack ),
    .X(_00478_));
 sky130_fd_sc_hd__nor2_1 _05814_ (.A(\u_semaphore.reg_ack ),
    .B(_01561_),
    .Y(_00476_));
 sky130_fd_sc_hd__o211a_1 _05815_ (.A1(net1329),
    .A2(_01544_),
    .B1(_01562_),
    .C1(\u_semaphore.reg_ack ),
    .X(_00477_));
 sky130_fd_sc_hd__and2_1 _05816_ (.A(net1243),
    .B(_01390_),
    .X(_01563_));
 sky130_fd_sc_hd__and3_1 _05817_ (.A(net1318),
    .B(\u_pwm.reg_ack_glbl ),
    .C(_01563_),
    .X(_00313_));
 sky130_fd_sc_hd__and3_1 _05818_ (.A(net1335),
    .B(\u_pwm.reg_ack_glbl ),
    .C(_01563_),
    .X(_00312_));
 sky130_fd_sc_hd__and4bb_1 _05819_ (.A_N(_01388_),
    .B_N(\u_pwm.reg_ack_glbl ),
    .C(net1255),
    .D(net1214),
    .X(_00311_));
 sky130_fd_sc_hd__nor2_1 _05820_ (.A(net1228),
    .B(_01532_),
    .Y(_01564_));
 sky130_fd_sc_hd__and2_1 _05821_ (.A(net1321),
    .B(_01564_),
    .X(_00354_));
 sky130_fd_sc_hd__and2_1 _05822_ (.A(net1327),
    .B(_01564_),
    .X(_00357_));
 sky130_fd_sc_hd__and2_1 _05823_ (.A(net1336),
    .B(_01564_),
    .X(_00356_));
 sky130_fd_sc_hd__nor2_2 _05824_ (.A(_00999_),
    .B(_01532_),
    .Y(_01565_));
 sky130_fd_sc_hd__and2_1 _05825_ (.A(net1321),
    .B(_01565_),
    .X(_00358_));
 sky130_fd_sc_hd__and2_1 _05826_ (.A(net1329),
    .B(_01565_),
    .X(_00361_));
 sky130_fd_sc_hd__and2_1 _05827_ (.A(net1336),
    .B(_01565_),
    .X(_00360_));
 sky130_fd_sc_hd__nor2_2 _05828_ (.A(_01115_),
    .B(_01532_),
    .Y(_01566_));
 sky130_fd_sc_hd__and2_1 _05829_ (.A(net1321),
    .B(_01566_),
    .X(_00362_));
 sky130_fd_sc_hd__and2_1 _05830_ (.A(net1327),
    .B(_01566_),
    .X(_00365_));
 sky130_fd_sc_hd__and2_1 _05831_ (.A(net1336),
    .B(_01566_),
    .X(_00364_));
 sky130_fd_sc_hd__and2_1 _05832_ (.A(net1321),
    .B(_01533_),
    .X(_00366_));
 sky130_fd_sc_hd__and2_1 _05833_ (.A(net1329),
    .B(_01533_),
    .X(_00369_));
 sky130_fd_sc_hd__and2_1 _05834_ (.A(net1336),
    .B(_01533_),
    .X(_00368_));
 sky130_fd_sc_hd__and4bb_1 _05835_ (.A_N(_01388_),
    .B_N(\u_pwm.reg_ack_pwm0 ),
    .C(net1255),
    .D(net1182),
    .X(_00352_));
 sky130_fd_sc_hd__and2_1 _05836_ (.A(net1313),
    .B(_01564_),
    .X(_00355_));
 sky130_fd_sc_hd__and2_1 _05837_ (.A(net1313),
    .B(_01565_),
    .X(_00359_));
 sky130_fd_sc_hd__and2_1 _05838_ (.A(net1313),
    .B(_01566_),
    .X(_00363_));
 sky130_fd_sc_hd__nor2_1 _05839_ (.A(net1222),
    .B(_01534_),
    .Y(_01567_));
 sky130_fd_sc_hd__and2_1 _05840_ (.A(net1318),
    .B(_01567_),
    .X(_00407_));
 sky130_fd_sc_hd__and2_1 _05841_ (.A(net1327),
    .B(_01567_),
    .X(_00410_));
 sky130_fd_sc_hd__and2_1 _05842_ (.A(net1335),
    .B(_01567_),
    .X(_00409_));
 sky130_fd_sc_hd__nor2_2 _05843_ (.A(_00999_),
    .B(_01534_),
    .Y(_01568_));
 sky130_fd_sc_hd__and2_1 _05844_ (.A(net1318),
    .B(_01568_),
    .X(_00411_));
 sky130_fd_sc_hd__and2_1 _05845_ (.A(net1328),
    .B(_01568_),
    .X(_00414_));
 sky130_fd_sc_hd__and2_1 _05846_ (.A(net1334),
    .B(_01568_),
    .X(_00413_));
 sky130_fd_sc_hd__nor2_2 _05847_ (.A(_01115_),
    .B(_01534_),
    .Y(_01569_));
 sky130_fd_sc_hd__and2_1 _05848_ (.A(net1318),
    .B(_01569_),
    .X(_00415_));
 sky130_fd_sc_hd__and2_1 _05849_ (.A(net1327),
    .B(_01569_),
    .X(_00418_));
 sky130_fd_sc_hd__and2_1 _05850_ (.A(net1334),
    .B(_01569_),
    .X(_00417_));
 sky130_fd_sc_hd__and2_1 _05851_ (.A(net1318),
    .B(_01535_),
    .X(_00419_));
 sky130_fd_sc_hd__and2_1 _05852_ (.A(net1327),
    .B(_01535_),
    .X(_00422_));
 sky130_fd_sc_hd__and2_1 _05853_ (.A(net1334),
    .B(_01535_),
    .X(_00421_));
 sky130_fd_sc_hd__and3b_1 _05854_ (.A_N(\u_pwm.reg_ack_pwm1 ),
    .B(_01118_),
    .C(_01389_),
    .X(_00405_));
 sky130_fd_sc_hd__and2_1 _05855_ (.A(net1311),
    .B(_01567_),
    .X(_00408_));
 sky130_fd_sc_hd__and2_1 _05856_ (.A(net1314),
    .B(_01568_),
    .X(_00412_));
 sky130_fd_sc_hd__and2_1 _05857_ (.A(net1311),
    .B(_01569_),
    .X(_00416_));
 sky130_fd_sc_hd__nor2_2 _05858_ (.A(net1221),
    .B(_01536_),
    .Y(_01570_));
 sky130_fd_sc_hd__and2_1 _05859_ (.A(net1318),
    .B(_01570_),
    .X(_00460_));
 sky130_fd_sc_hd__and2_1 _05860_ (.A(net1326),
    .B(_01570_),
    .X(_00463_));
 sky130_fd_sc_hd__and2_1 _05861_ (.A(net1333),
    .B(_01570_),
    .X(_00462_));
 sky130_fd_sc_hd__nor2_4 _05862_ (.A(_00999_),
    .B(_01536_),
    .Y(_01571_));
 sky130_fd_sc_hd__and2_1 _05863_ (.A(net1318),
    .B(_01571_),
    .X(_00464_));
 sky130_fd_sc_hd__and2_1 _05864_ (.A(net1326),
    .B(_01571_),
    .X(_00467_));
 sky130_fd_sc_hd__and2_1 _05865_ (.A(net1333),
    .B(_01571_),
    .X(_00466_));
 sky130_fd_sc_hd__nor2_4 _05866_ (.A(_01115_),
    .B(_01536_),
    .Y(_01572_));
 sky130_fd_sc_hd__and2_1 _05867_ (.A(net62),
    .B(_01572_),
    .X(_00468_));
 sky130_fd_sc_hd__and2_1 _05868_ (.A(net1326),
    .B(_01572_),
    .X(_00471_));
 sky130_fd_sc_hd__and2_1 _05869_ (.A(net1333),
    .B(_01572_),
    .X(_00470_));
 sky130_fd_sc_hd__and2_1 _05870_ (.A(net62),
    .B(_01537_),
    .X(_00472_));
 sky130_fd_sc_hd__and2_1 _05871_ (.A(net1326),
    .B(_01537_),
    .X(_00475_));
 sky130_fd_sc_hd__and2_1 _05872_ (.A(net1333),
    .B(_01537_),
    .X(_00474_));
 sky130_fd_sc_hd__nor3_2 _05873_ (.A(\u_pwm.reg_ack_pwm2 ),
    .B(_01145_),
    .C(_01388_),
    .Y(_00458_));
 sky130_fd_sc_hd__and2_1 _05874_ (.A(net1310),
    .B(_01570_),
    .X(_00461_));
 sky130_fd_sc_hd__and2_1 _05875_ (.A(net1310),
    .B(_01571_),
    .X(_00465_));
 sky130_fd_sc_hd__and2_1 _05876_ (.A(net1310),
    .B(_01572_),
    .X(_00469_));
 sky130_fd_sc_hd__nand2b_1 _05877_ (.A_N(net1388),
    .B(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .Y(net503));
 sky130_fd_sc_hd__and2b_1 _05878_ (.A_N(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .B(\u_gpio.cfg_gpio_dir_sel[21] ),
    .X(_01573_));
 sky130_fd_sc_hd__a22o_2 _05879_ (.A1(net1377),
    .A2(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .B1(_01573_),
    .B2(\u_gpio.cfg_gpio_out_data[21] ),
    .X(net310));
 sky130_fd_sc_hd__and2b_1 _05880_ (.A_N(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .B(\u_gpio.cfg_gpio_dir_sel[20] ),
    .X(_01574_));
 sky130_fd_sc_hd__a22o_2 _05881_ (.A1(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .A2(net42),
    .B1(_01574_),
    .B2(\u_gpio.cfg_gpio_out_data[20] ),
    .X(net309));
 sky130_fd_sc_hd__and2_1 _05882_ (.A(\u_gpio.cfg_gpio_out_data[19] ),
    .B(\u_gpio.cfg_gpio_dir_sel[19] ),
    .X(_01575_));
 sky130_fd_sc_hd__a31o_2 _05883_ (.A1(net1399),
    .A2(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .A3(_00935_),
    .B1(_01575_),
    .X(net308));
 sky130_fd_sc_hd__and2_1 _05884_ (.A(\u_gpio.cfg_gpio_out_data[18] ),
    .B(\u_gpio.cfg_gpio_dir_sel[18] ),
    .X(_01576_));
 sky130_fd_sc_hd__mux2_2 _05885_ (.A0(_01576_),
    .A1(net195),
    .S(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .X(net307));
 sky130_fd_sc_hd__nor2_2 _05886_ (.A(\u_gpio.cfg_gpio_dir_sel[13] ),
    .B(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .Y(net266));
 sky130_fd_sc_hd__and2_1 _05887_ (.A(\u_gpio.cfg_gpio_out_data[13] ),
    .B(\u_gpio.cfg_gpio_dir_sel[13] ),
    .X(_01577_));
 sky130_fd_sc_hd__mux2_2 _05888_ (.A0(_01577_),
    .A1(net153),
    .S(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .X(net304));
 sky130_fd_sc_hd__and2_1 _05889_ (.A(\u_gpio.cfg_gpio_out_data[12] ),
    .B(\u_gpio.cfg_gpio_dir_sel[12] ),
    .X(_01578_));
 sky130_fd_sc_hd__mux2_1 _05890_ (.A0(_01578_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[12] ),
    .X(_01579_));
 sky130_fd_sc_hd__mux2_2 _05891_ (.A0(_01579_),
    .A1(net152),
    .S(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .X(net303));
 sky130_fd_sc_hd__or2_4 _05892_ (.A(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .B(net34),
    .X(net463));
 sky130_fd_sc_hd__or3b_1 _05893_ (.A(\u_gpio.cfg_gpio_dir_sel[11] ),
    .B(net463),
    .C_N(net158),
    .X(_01580_));
 sky130_fd_sc_hd__a21bo_1 _05894_ (.A1(\u_gpio.cfg_gpio_out_data[11] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[11] ),
    .B1_N(_01580_),
    .X(_01581_));
 sky130_fd_sc_hd__mux2_1 _05895_ (.A0(_01581_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[11] ),
    .X(_01582_));
 sky130_fd_sc_hd__xor2_2 _05896_ (.A(\u_pwm.u_pwm_2.cfg_pwm_inv ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_wfm_r ),
    .X(_01583_));
 sky130_fd_sc_hd__mux2_2 _05897_ (.A0(_01582_),
    .A1(_01583_),
    .S(\u_glbl_reg.cfg_multi_func_sel[5] ),
    .X(net301));
 sky130_fd_sc_hd__xor2_2 _05898_ (.A(\u_pwm.u_pwm_1.cfg_pwm_inv ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_wfm_r ),
    .X(_01584_));
 sky130_fd_sc_hd__and3b_1 _05899_ (.A_N(\u_gpio.cfg_gpio_out_type[10] ),
    .B(\u_gpio.cfg_gpio_dir_sel[10] ),
    .C(\u_gpio.cfg_gpio_out_data[10] ),
    .X(_01585_));
 sky130_fd_sc_hd__a21o_1 _05900_ (.A1(net1078),
    .A2(\u_gpio.cfg_gpio_out_type[10] ),
    .B1(_01585_),
    .X(_01586_));
 sky130_fd_sc_hd__mux2_1 _05901_ (.A0(_01586_),
    .A1(net154),
    .S(\u_glbl_reg.cfg_multi_func_sel[11] ),
    .X(_01587_));
 sky130_fd_sc_hd__mux2_2 _05902_ (.A0(_01587_),
    .A1(_01584_),
    .S(\u_glbl_reg.cfg_multi_func_sel[4] ),
    .X(net300));
 sky130_fd_sc_hd__xor2_4 _05903_ (.A(\u_pwm.u_pwm_0.cfg_pwm_inv ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_wfm_r ),
    .X(_01588_));
 sky130_fd_sc_hd__and3b_1 _05904_ (.A_N(\u_gpio.cfg_gpio_out_type[9] ),
    .B(\u_gpio.cfg_gpio_dir_sel[9] ),
    .C(\u_gpio.cfg_gpio_out_data[9] ),
    .X(_01589_));
 sky130_fd_sc_hd__a21o_1 _05905_ (.A1(net1078),
    .A2(\u_gpio.cfg_gpio_out_type[9] ),
    .B1(_01589_),
    .X(_01590_));
 sky130_fd_sc_hd__mux2_1 _05906_ (.A0(_01590_),
    .A1(net155),
    .S(\u_glbl_reg.cfg_multi_func_sel[12] ),
    .X(_01591_));
 sky130_fd_sc_hd__mux2_2 _05907_ (.A0(_01591_),
    .A1(_01588_),
    .S(\u_glbl_reg.cfg_multi_func_sel[3] ),
    .X(net299));
 sky130_fd_sc_hd__and2_1 _05908_ (.A(\u_gpio.cfg_gpio_out_data[8] ),
    .B(\u_gpio.cfg_gpio_dir_sel[8] ),
    .X(_01592_));
 sky130_fd_sc_hd__mux2_1 _05909_ (.A0(_01592_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[8] ),
    .X(net298));
 sky130_fd_sc_hd__and2_1 _05910_ (.A(\u_gpio.cfg_gpio_out_data[31] ),
    .B(\u_gpio.cfg_gpio_dir_sel[31] ),
    .X(_01593_));
 sky130_fd_sc_hd__mux2_1 _05911_ (.A0(_01593_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[31] ),
    .X(_01594_));
 sky130_fd_sc_hd__mux2_2 _05912_ (.A0(net564),
    .A1(net47),
    .S(\u_glbl_reg.cfg_multi_func_sel[17] ),
    .X(net297));
 sky130_fd_sc_hd__and2_1 _05913_ (.A(\u_gpio.cfg_gpio_out_data[30] ),
    .B(\u_gpio.cfg_gpio_dir_sel[30] ),
    .X(_01595_));
 sky130_fd_sc_hd__mux2_1 _05914_ (.A0(_01595_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[30] ),
    .X(_01596_));
 sky130_fd_sc_hd__mux2_1 _05915_ (.A0(_01596_),
    .A1(net156),
    .S(\u_glbl_reg.cfg_multi_func_sel[13] ),
    .X(_01597_));
 sky130_fd_sc_hd__mux2_1 _05916_ (.A0(_01597_),
    .A1(_01583_),
    .S(\u_glbl_reg.cfg_multi_func_sel[2] ),
    .X(net296));
 sky130_fd_sc_hd__and2_1 _05917_ (.A(\u_gpio.cfg_gpio_out_data[29] ),
    .B(\u_gpio.cfg_gpio_dir_sel[29] ),
    .X(_01598_));
 sky130_fd_sc_hd__mux2_1 _05918_ (.A0(_01598_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[29] ),
    .X(_01599_));
 sky130_fd_sc_hd__mux2_1 _05919_ (.A0(_01599_),
    .A1(net157),
    .S(\u_glbl_reg.cfg_multi_func_sel[14] ),
    .X(_01600_));
 sky130_fd_sc_hd__mux2_4 _05920_ (.A0(_01600_),
    .A1(_01584_),
    .S(\u_glbl_reg.cfg_multi_func_sel[1] ),
    .X(net295));
 sky130_fd_sc_hd__nor2_4 _05921_ (.A(\u_gpio.cfg_gpio_dir_sel[15] ),
    .B(\u_gpio.cfg_gpio_out_type[15] ),
    .Y(net256));
 sky130_fd_sc_hd__and2_1 _05922_ (.A(\u_gpio.cfg_gpio_out_data[15] ),
    .B(\u_gpio.cfg_gpio_dir_sel[15] ),
    .X(_01601_));
 sky130_fd_sc_hd__mux2_4 _05923_ (.A0(_01601_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[15] ),
    .X(net294));
 sky130_fd_sc_hd__nor2_4 _05924_ (.A(\u_gpio.cfg_gpio_dir_sel[14] ),
    .B(\u_gpio.cfg_gpio_out_type[14] ),
    .Y(net255));
 sky130_fd_sc_hd__and2_1 _05925_ (.A(\u_gpio.cfg_gpio_out_data[14] ),
    .B(\u_gpio.cfg_gpio_dir_sel[14] ),
    .X(_01602_));
 sky130_fd_sc_hd__mux2_4 _05926_ (.A0(_01602_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[14] ),
    .X(net293));
 sky130_fd_sc_hd__and2_1 _05927_ (.A(\u_gpio.cfg_gpio_out_data[28] ),
    .B(\u_gpio.cfg_gpio_dir_sel[28] ),
    .X(_01603_));
 sky130_fd_sc_hd__mux2_1 _05928_ (.A0(_01603_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[28] ),
    .X(_01604_));
 sky130_fd_sc_hd__mux2_4 _05929_ (.A0(_01604_),
    .A1(net192),
    .S(\u_glbl_reg.cfg_multi_func_sel[9] ),
    .X(net292));
 sky130_fd_sc_hd__and2_1 _05930_ (.A(\u_gpio.cfg_gpio_out_data[27] ),
    .B(\u_gpio.cfg_gpio_dir_sel[27] ),
    .X(_01605_));
 sky130_fd_sc_hd__mux2_1 _05931_ (.A0(_01605_),
    .A1(net1078),
    .S(\u_gpio.cfg_gpio_out_type[27] ),
    .X(_01606_));
 sky130_fd_sc_hd__mux2_4 _05932_ (.A0(_01606_),
    .A1(_01588_),
    .S(\u_glbl_reg.cfg_multi_func_sel[0] ),
    .X(net328));
 sky130_fd_sc_hd__and2_1 _05933_ (.A(\u_gpio.cfg_gpio_out_data[26] ),
    .B(\u_gpio.cfg_gpio_dir_sel[26] ),
    .X(_01607_));
 sky130_fd_sc_hd__mux2_4 _05934_ (.A0(_01607_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[26] ),
    .X(net327));
 sky130_fd_sc_hd__and3b_1 _05935_ (.A_N(\u_gpio.cfg_gpio_out_type[25] ),
    .B(\u_gpio.cfg_gpio_dir_sel[25] ),
    .C(\u_gpio.cfg_gpio_out_data[25] ),
    .X(_01608_));
 sky130_fd_sc_hd__a21o_1 _05936_ (.A1(net1079),
    .A2(\u_gpio.cfg_gpio_out_type[25] ),
    .B1(_01608_),
    .X(_01609_));
 sky130_fd_sc_hd__mux2_1 _05937_ (.A0(_01609_),
    .A1(net191),
    .S(\u_glbl_reg.cfg_multi_func_sel[8] ),
    .X(_01610_));
 sky130_fd_sc_hd__mux2_2 _05938_ (.A0(_01610_),
    .A1(net193),
    .S(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .X(net326));
 sky130_fd_sc_hd__nor2_1 _05939_ (.A(\u_gpio.cfg_gpio_dir_sel[24] ),
    .B(\u_gpio.cfg_gpio_out_type[24] ),
    .Y(_01611_));
 sky130_fd_sc_hd__and2_1 _05940_ (.A(\u_gpio.cfg_gpio_out_data[24] ),
    .B(\u_gpio.cfg_gpio_dir_sel[24] ),
    .X(_01612_));
 sky130_fd_sc_hd__mux2_4 _05941_ (.A0(_01612_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[24] ),
    .X(net325));
 sky130_fd_sc_hd__nor2_4 _05942_ (.A(\u_gpio.cfg_gpio_dir_sel[22] ),
    .B(\u_gpio.cfg_gpio_out_type[22] ),
    .Y(net286));
 sky130_fd_sc_hd__and2_1 _05943_ (.A(\u_gpio.cfg_gpio_out_data[22] ),
    .B(\u_gpio.cfg_gpio_dir_sel[22] ),
    .X(_01613_));
 sky130_fd_sc_hd__mux2_4 _05944_ (.A0(_01613_),
    .A1(net1079),
    .S(\u_gpio.cfg_gpio_out_type[22] ),
    .X(net324));
 sky130_fd_sc_hd__mux2_2 _05945_ (.A0(_00937_),
    .A1(net1414),
    .S(net1109),
    .X(net285));
 sky130_fd_sc_hd__a21oi_4 _05946_ (.A1(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .A2(_00938_),
    .B1(_01573_),
    .Y(net272));
 sky130_fd_sc_hd__a21oi_4 _05947_ (.A1(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .A2(_00939_),
    .B1(_01574_),
    .Y(net271));
 sky130_fd_sc_hd__mux2_2 _05948_ (.A0(_00935_),
    .A1(net1398),
    .S(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .X(net270));
 sky130_fd_sc_hd__mux2_2 _05949_ (.A0(_00936_),
    .A1(net1398),
    .S(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .X(net269));
 sky130_fd_sc_hd__nor3_4 _05950_ (.A(\u_gpio.cfg_gpio_dir_sel[28] ),
    .B(\u_gpio.cfg_gpio_out_type[28] ),
    .C(\u_glbl_reg.cfg_multi_func_sel[9] ),
    .Y(net254));
 sky130_fd_sc_hd__o21ba_1 _05951_ (.A1(\u_gpio.cfg_gpio_dir_sel[27] ),
    .A2(\u_gpio.cfg_gpio_out_type[27] ),
    .B1_N(\u_glbl_reg.cfg_multi_func_sel[7] ),
    .X(_01614_));
 sky130_fd_sc_hd__nor2_4 _05952_ (.A(\u_glbl_reg.cfg_multi_func_sel[0] ),
    .B(_01614_),
    .Y(net290));
 sky130_fd_sc_hd__nor4_4 _05953_ (.A(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .B(\u_gpio.cfg_gpio_dir_sel[25] ),
    .C(\u_gpio.cfg_gpio_out_type[25] ),
    .D(\u_glbl_reg.cfg_multi_func_sel[8] ),
    .Y(net288));
 sky130_fd_sc_hd__or2_1 _05954_ (.A(net1400),
    .B(net463),
    .X(net462));
 sky130_fd_sc_hd__nand2b_4 _05955_ (.A_N(net19),
    .B(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .Y(net506));
 sky130_fd_sc_hd__nand2b_1 _05956_ (.A_N(net20),
    .B(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .Y(net505));
 sky130_fd_sc_hd__nand2b_4 _05957_ (.A_N(net1392),
    .B(net1109),
    .Y(net453));
 sky130_fd_sc_hd__mux2_2 _05958_ (.A0(\u_gpio.cfg_gpio_out_data[0] ),
    .A1(net1405),
    .S(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .X(net291));
 sky130_fd_sc_hd__mux2_2 _05959_ (.A0(\u_gpio.cfg_gpio_out_data[1] ),
    .A1(net1404),
    .S(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .X(net302));
 sky130_fd_sc_hd__mux2_2 _05960_ (.A0(\u_gpio.cfg_gpio_out_data[2] ),
    .A1(net1402),
    .S(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .X(net313));
 sky130_fd_sc_hd__mux2_2 _05961_ (.A0(\u_gpio.cfg_gpio_out_data[3] ),
    .A1(net1401),
    .S(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .X(net322));
 sky130_fd_sc_hd__mux2_2 _05962_ (.A0(\u_gpio.cfg_gpio_out_data[4] ),
    .A1(net1415),
    .S(net1109),
    .X(net323));
 sky130_fd_sc_hd__xnor2_1 _05963_ (.A(\u_glbl_reg.u_dbgclk.high_count[1] ),
    .B(\u_glbl_reg.u_dbgclk.high_count[0] ),
    .Y(_00040_));
 sky130_fd_sc_hd__o21ai_1 _05964_ (.A1(\u_glbl_reg.u_dbgclk.high_count[1] ),
    .A2(\u_glbl_reg.u_dbgclk.high_count[0] ),
    .B1(\u_glbl_reg.u_dbgclk.high_count[2] ),
    .Y(_01615_));
 sky130_fd_sc_hd__nand2_1 _05965_ (.A(_01106_),
    .B(_01615_),
    .Y(_00041_));
 sky130_fd_sc_hd__and2_1 _05966_ (.A(\u_glbl_reg.u_dbgclk.high_count[3] ),
    .B(_01106_),
    .X(_00042_));
 sky130_fd_sc_hd__and2b_1 _05967_ (.A_N(\u_glbl_reg.u_dbgclk.low_count[0] ),
    .B(_01108_),
    .X(_00046_));
 sky130_fd_sc_hd__o21ba_1 _05968_ (.A1(\u_glbl_reg.u_dbgclk.low_count[3] ),
    .A2(\u_glbl_reg.u_dbgclk.low_count[2] ),
    .B1_N(_01107_),
    .X(_01616_));
 sky130_fd_sc_hd__a21o_1 _05969_ (.A1(\u_glbl_reg.u_dbgclk.low_count[0] ),
    .A2(\u_glbl_reg.u_dbgclk.low_count[1] ),
    .B1(_01616_),
    .X(_00047_));
 sky130_fd_sc_hd__mux2_1 _05970_ (.A0(_01616_),
    .A1(_01107_),
    .S(\u_glbl_reg.u_dbgclk.low_count[2] ),
    .X(_00048_));
 sky130_fd_sc_hd__o21ai_1 _05971_ (.A1(\u_glbl_reg.u_dbgclk.low_count[2] ),
    .A2(_01107_),
    .B1(\u_glbl_reg.u_dbgclk.low_count[3] ),
    .Y(_01617_));
 sky130_fd_sc_hd__nand2_1 _05972_ (.A(_01108_),
    .B(_01617_),
    .Y(_00049_));
 sky130_fd_sc_hd__xnor2_1 _05973_ (.A(\u_glbl_reg.cfg_ref_pll_div[0] ),
    .B(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .Y(_01618_));
 sky130_fd_sc_hd__a21oi_1 _05974_ (.A1(_00055_),
    .A2(_01618_),
    .B1(\u_glbl_reg.u_pll_ref_clk.high_count[0] ),
    .Y(_00050_));
 sky130_fd_sc_hd__nand2_1 _05975_ (.A(\u_glbl_reg.u_pll_ref_clk.high_count[1] ),
    .B(\u_glbl_reg.u_pll_ref_clk.high_count[0] ),
    .Y(_01619_));
 sky130_fd_sc_hd__a21oi_1 _05976_ (.A1(\u_glbl_reg.cfg_ref_pll_div[0] ),
    .A2(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .B1(\u_glbl_reg.cfg_ref_pll_div[2] ),
    .Y(_01620_));
 sky130_fd_sc_hd__and3_1 _05977_ (.A(\u_glbl_reg.cfg_ref_pll_div[0] ),
    .B(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .C(\u_glbl_reg.cfg_ref_pll_div[2] ),
    .X(_01621_));
 sky130_fd_sc_hd__o21ba_1 _05978_ (.A1(_01620_),
    .A2(_01621_),
    .B1_N(\u_glbl_reg.u_pll_ref_clk.high_count[2] ),
    .X(_01622_));
 sky130_fd_sc_hd__o21ai_1 _05979_ (.A1(_01109_),
    .A2(_01622_),
    .B1(_01619_),
    .Y(_00051_));
 sky130_fd_sc_hd__and2_1 _05980_ (.A(\u_glbl_reg.u_pll_ref_clk.high_count[2] ),
    .B(_01109_),
    .X(_01623_));
 sky130_fd_sc_hd__a21o_1 _05981_ (.A1(_00055_),
    .A2(_01621_),
    .B1(_01623_),
    .X(_00052_));
 sky130_fd_sc_hd__a21oi_1 _05982_ (.A1(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .A2(_01111_),
    .B1(\u_glbl_reg.u_pll_ref_clk.low_count[0] ),
    .Y(_00056_));
 sky130_fd_sc_hd__xor2_1 _05983_ (.A(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .B(\u_glbl_reg.cfg_ref_pll_div[2] ),
    .X(_01624_));
 sky130_fd_sc_hd__o21ba_1 _05984_ (.A1(\u_glbl_reg.u_pll_ref_clk.low_count[2] ),
    .A2(_01624_),
    .B1_N(_01110_),
    .X(_01625_));
 sky130_fd_sc_hd__a21o_1 _05985_ (.A1(\u_glbl_reg.u_pll_ref_clk.low_count[0] ),
    .A2(\u_glbl_reg.u_pll_ref_clk.low_count[1] ),
    .B1(_01625_),
    .X(_00057_));
 sky130_fd_sc_hd__and2_1 _05986_ (.A(\u_glbl_reg.u_pll_ref_clk.low_count[2] ),
    .B(_01110_),
    .X(_01626_));
 sky130_fd_sc_hd__a31o_1 _05987_ (.A1(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .A2(\u_glbl_reg.cfg_ref_pll_div[2] ),
    .A3(_01111_),
    .B1(_01626_),
    .X(_00058_));
 sky130_fd_sc_hd__mux2_1 _05988_ (.A0(net1427),
    .A1(net162),
    .S(net1205),
    .X(_00121_));
 sky130_fd_sc_hd__and2b_1 _05989_ (.A_N(net1205),
    .B(net1418),
    .X(_00122_));
 sky130_fd_sc_hd__and2b_1 _05990_ (.A_N(net1204),
    .B(net1288),
    .X(_00092_));
 sky130_fd_sc_hd__and2b_1 _05991_ (.A_N(net1203),
    .B(net1644),
    .X(_00093_));
 sky130_fd_sc_hd__and2b_1 _05992_ (.A_N(net1205),
    .B(net1638),
    .X(_00094_));
 sky130_fd_sc_hd__and2b_1 _05993_ (.A_N(net1204),
    .B(net1628),
    .X(_00095_));
 sky130_fd_sc_hd__and2b_1 _05994_ (.A_N(net1204),
    .B(net1621),
    .X(_00096_));
 sky130_fd_sc_hd__and2b_1 _05995_ (.A_N(net1204),
    .B(net1615),
    .X(_00097_));
 sky130_fd_sc_hd__and2b_1 _05996_ (.A_N(net1203),
    .B(net1603),
    .X(_00098_));
 sky130_fd_sc_hd__and2b_1 _05997_ (.A_N(net1203),
    .B(net1595),
    .X(_00099_));
 sky130_fd_sc_hd__and2b_1 _05998_ (.A_N(net1203),
    .B(net1586),
    .X(_00100_));
 sky130_fd_sc_hd__and2b_1 _05999_ (.A_N(net1204),
    .B(net1579),
    .X(_00101_));
 sky130_fd_sc_hd__and2b_1 _06000_ (.A_N(net1203),
    .B(net1564),
    .X(_00103_));
 sky130_fd_sc_hd__and2b_1 _06001_ (.A_N(net1203),
    .B(net1556),
    .X(_00104_));
 sky130_fd_sc_hd__and2b_1 _06002_ (.A_N(net1203),
    .B(net1549),
    .X(_00105_));
 sky130_fd_sc_hd__and2b_1 _06003_ (.A_N(net1203),
    .B(net1541),
    .X(_00106_));
 sky130_fd_sc_hd__and2b_1 _06004_ (.A_N(net1202),
    .B(net1535),
    .X(_00107_));
 sky130_fd_sc_hd__and2b_1 _06005_ (.A_N(net1202),
    .B(net1526),
    .X(_00108_));
 sky130_fd_sc_hd__and2b_1 _06006_ (.A_N(net1201),
    .B(net1519),
    .X(_00109_));
 sky130_fd_sc_hd__and2b_1 _06007_ (.A_N(net1201),
    .B(net1512),
    .X(_00110_));
 sky130_fd_sc_hd__and2b_1 _06008_ (.A_N(net1202),
    .B(net1505),
    .X(_00111_));
 sky130_fd_sc_hd__and2b_1 _06009_ (.A_N(net1201),
    .B(net1498),
    .X(_00112_));
 sky130_fd_sc_hd__and2b_1 _06010_ (.A_N(net1202),
    .B(net1481),
    .X(_00114_));
 sky130_fd_sc_hd__and2b_1 _06011_ (.A_N(net1202),
    .B(net1474),
    .X(_00115_));
 sky130_fd_sc_hd__and2_1 _06012_ (.A(_00795_),
    .B(net164),
    .X(_01627_));
 sky130_fd_sc_hd__a21o_1 _06013_ (.A1(net1603),
    .A2(net774),
    .B1(_01627_),
    .X(_00032_));
 sky130_fd_sc_hd__a21o_1 _06014_ (.A1(net1595),
    .A2(net774),
    .B1(_01627_),
    .X(_00033_));
 sky130_fd_sc_hd__a21o_1 _06015_ (.A1(net1586),
    .A2(net774),
    .B1(_01627_),
    .X(_00034_));
 sky130_fd_sc_hd__a21o_1 _06016_ (.A1(net1579),
    .A2(net774),
    .B1(_01627_),
    .X(_00035_));
 sky130_fd_sc_hd__mux2_1 _06017_ (.A0(net163),
    .A1(net1519),
    .S(net735),
    .X(_00036_));
 sky130_fd_sc_hd__mux2_1 _06018_ (.A0(net163),
    .A1(net1512),
    .S(net735),
    .X(_00037_));
 sky130_fd_sc_hd__xnor2_1 _06019_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ),
    .B(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .Y(_01628_));
 sky130_fd_sc_hd__a21oi_1 _06020_ (.A1(_00194_),
    .A2(_01628_),
    .B1(\u_glbl_reg.u_rtcclk.high_count[0] ),
    .Y(_00187_));
 sky130_fd_sc_hd__nand2_1 _06021_ (.A(\u_glbl_reg.u_rtcclk.high_count[0] ),
    .B(\u_glbl_reg.u_rtcclk.high_count[1] ),
    .Y(_01629_));
 sky130_fd_sc_hd__a21oi_1 _06022_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ),
    .A2(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .B1(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .Y(_01630_));
 sky130_fd_sc_hd__and3_1 _06023_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ),
    .B(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .C(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .X(_01631_));
 sky130_fd_sc_hd__o21a_1 _06024_ (.A1(_01630_),
    .A2(_01631_),
    .B1(_00194_),
    .X(_01632_));
 sky130_fd_sc_hd__a21oi_1 _06025_ (.A1(_01135_),
    .A2(_01629_),
    .B1(_01632_),
    .Y(_00188_));
 sky130_fd_sc_hd__nand2_1 _06026_ (.A(\u_glbl_reg.u_rtcclk.high_count[2] ),
    .B(_01135_),
    .Y(_01633_));
 sky130_fd_sc_hd__and3_1 _06027_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .B(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .C(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ),
    .X(_01634_));
 sky130_fd_sc_hd__and2_1 _06028_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ),
    .B(_01634_),
    .X(_01635_));
 sky130_fd_sc_hd__nor2_1 _06029_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ),
    .B(_01631_),
    .Y(_01636_));
 sky130_fd_sc_hd__o21a_1 _06030_ (.A1(_01635_),
    .A2(_01636_),
    .B1(_00194_),
    .X(_01637_));
 sky130_fd_sc_hd__a21oi_1 _06031_ (.A1(_01136_),
    .A2(_01633_),
    .B1(_01637_),
    .Y(_00189_));
 sky130_fd_sc_hd__nand2_1 _06032_ (.A(\u_glbl_reg.u_rtcclk.high_count[3] ),
    .B(_01136_),
    .Y(_01638_));
 sky130_fd_sc_hd__nor2_1 _06033_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ),
    .B(_01635_),
    .Y(_01639_));
 sky130_fd_sc_hd__and3_1 _06034_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ),
    .B(_00194_),
    .C(_01635_),
    .X(_01640_));
 sky130_fd_sc_hd__a221oi_1 _06035_ (.A1(_01137_),
    .A2(_01638_),
    .B1(_01639_),
    .B2(_00194_),
    .C1(_01640_),
    .Y(_00190_));
 sky130_fd_sc_hd__a21o_1 _06036_ (.A1(\u_glbl_reg.u_rtcclk.high_count[4] ),
    .A2(_01137_),
    .B1(_01640_),
    .X(_00191_));
 sky130_fd_sc_hd__a21oi_1 _06037_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .A2(_01142_),
    .B1(\u_glbl_reg.u_rtcclk.low_count[0] ),
    .Y(_00195_));
 sky130_fd_sc_hd__and2_1 _06038_ (.A(\u_glbl_reg.u_rtcclk.low_count[1] ),
    .B(\u_glbl_reg.u_rtcclk.low_count[0] ),
    .X(_01641_));
 sky130_fd_sc_hd__xor2_1 _06039_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .B(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .X(_01642_));
 sky130_fd_sc_hd__o22a_1 _06040_ (.A1(_01138_),
    .A2(_01641_),
    .B1(_01642_),
    .B2(_01143_),
    .X(_00196_));
 sky130_fd_sc_hd__o21ai_1 _06041_ (.A1(\u_glbl_reg.u_rtcclk.low_count[1] ),
    .A2(\u_glbl_reg.u_rtcclk.low_count[0] ),
    .B1(\u_glbl_reg.u_rtcclk.low_count[2] ),
    .Y(_01643_));
 sky130_fd_sc_hd__a21oi_1 _06042_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .A2(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .B1(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ),
    .Y(_01644_));
 sky130_fd_sc_hd__nor2_1 _06043_ (.A(_01634_),
    .B(_01644_),
    .Y(_01645_));
 sky130_fd_sc_hd__o2bb2a_1 _06044_ (.A1_N(_01139_),
    .A2_N(_01643_),
    .B1(_01645_),
    .B2(_01143_),
    .X(_00197_));
 sky130_fd_sc_hd__and2_1 _06045_ (.A(\u_glbl_reg.u_rtcclk.low_count[3] ),
    .B(_01139_),
    .X(_01646_));
 sky130_fd_sc_hd__xor2_1 _06046_ (.A(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ),
    .B(_01634_),
    .X(_01647_));
 sky130_fd_sc_hd__o22a_1 _06047_ (.A1(_01141_),
    .A2(_01646_),
    .B1(_01647_),
    .B2(_01143_),
    .X(_00198_));
 sky130_fd_sc_hd__and2_1 _06048_ (.A(\u_glbl_reg.u_rtcclk.low_count[4] ),
    .B(_01140_),
    .X(_01648_));
 sky130_fd_sc_hd__a31o_1 _06049_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ),
    .A2(_01142_),
    .A3(_01634_),
    .B1(_01648_),
    .X(_00199_));
 sky130_fd_sc_hd__nor2_1 _06050_ (.A(net1055),
    .B(\u_glbl_reg.reg_12[15] ),
    .Y(_01649_));
 sky130_fd_sc_hd__or2_1 _06051_ (.A(net1055),
    .B(\u_glbl_reg.reg_12[15] ),
    .X(_01650_));
 sky130_fd_sc_hd__a22o_1 _06052_ (.A1(net1534),
    .A2(net1045),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net598),
    .X(_00216_));
 sky130_fd_sc_hd__a22o_1 _06053_ (.A1(net1526),
    .A2(net1044),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00217_));
 sky130_fd_sc_hd__a22o_1 _06054_ (.A1(net1519),
    .A2(net1045),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net598),
    .X(_00218_));
 sky130_fd_sc_hd__a22o_1 _06055_ (.A1(net1512),
    .A2(net1044),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00219_));
 sky130_fd_sc_hd__a22o_1 _06056_ (.A1(net1505),
    .A2(net1045),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net598),
    .X(_00220_));
 sky130_fd_sc_hd__a22o_1 _06057_ (.A1(net1498),
    .A2(net1044),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00221_));
 sky130_fd_sc_hd__and2_1 _06058_ (.A(net1481),
    .B(net1045),
    .X(_00223_));
 sky130_fd_sc_hd__a22o_1 _06059_ (.A1(net1293),
    .A2(net1046),
    .B1(\u_glbl_reg.reg_12[0] ),
    .B2(net599),
    .X(_00200_));
 sky130_fd_sc_hd__a22o_1 _06060_ (.A1(net1572),
    .A2(net1047),
    .B1(\u_glbl_reg.reg_12[1] ),
    .B2(net599),
    .X(_00211_));
 sky130_fd_sc_hd__a22o_1 _06061_ (.A1(net1488),
    .A2(net1046),
    .B1(\u_glbl_reg.reg_12[2] ),
    .B2(net599),
    .X(_00222_));
 sky130_fd_sc_hd__a22o_1 _06062_ (.A1(net1466),
    .A2(net1047),
    .B1(\u_glbl_reg.reg_12[3] ),
    .B2(net599),
    .X(_00225_));
 sky130_fd_sc_hd__a22o_1 _06063_ (.A1(net1457),
    .A2(net1046),
    .B1(\u_glbl_reg.reg_12[0] ),
    .B2(net599),
    .X(_00226_));
 sky130_fd_sc_hd__a22o_1 _06064_ (.A1(net1448),
    .A2(net1047),
    .B1(\u_glbl_reg.reg_12[1] ),
    .B2(net599),
    .X(_00227_));
 sky130_fd_sc_hd__a22o_1 _06065_ (.A1(net1441),
    .A2(net1046),
    .B1(\u_glbl_reg.reg_12[2] ),
    .B2(net599),
    .X(_00228_));
 sky130_fd_sc_hd__a22o_1 _06066_ (.A1(net1433),
    .A2(net1047),
    .B1(\u_glbl_reg.reg_12[3] ),
    .B2(net599),
    .X(_00229_));
 sky130_fd_sc_hd__a22o_1 _06067_ (.A1(net1427),
    .A2(net1055),
    .B1(\u_glbl_reg.reg_12[4] ),
    .B2(net600),
    .X(_00230_));
 sky130_fd_sc_hd__o22a_1 _06068_ (.A1(net1419),
    .A2(_00796_),
    .B1(\u_glbl_reg.reg_12[5] ),
    .B2(_01650_),
    .X(_00231_));
 sky130_fd_sc_hd__a22o_1 _06069_ (.A1(net1286),
    .A2(net1055),
    .B1(\u_glbl_reg.reg_12[6] ),
    .B2(net600),
    .X(_00201_));
 sky130_fd_sc_hd__o22a_1 _06070_ (.A1(net1644),
    .A2(_00796_),
    .B1(\u_glbl_reg.reg_12[7] ),
    .B2(_01650_),
    .X(_00202_));
 sky130_fd_sc_hd__o22a_1 _06071_ (.A1(net1638),
    .A2(_00796_),
    .B1(\u_glbl_reg.reg_12[8] ),
    .B2(_01650_),
    .X(_00203_));
 sky130_fd_sc_hd__o22a_1 _06072_ (.A1(net1630),
    .A2(_00796_),
    .B1(\u_glbl_reg.reg_12[9] ),
    .B2(_01650_),
    .X(_00204_));
 sky130_fd_sc_hd__a22o_1 _06073_ (.A1(net1623),
    .A2(net1055),
    .B1(\u_glbl_reg.reg_12[10] ),
    .B2(net600),
    .X(_00205_));
 sky130_fd_sc_hd__and2_1 _06074_ (.A(net1613),
    .B(net1055),
    .X(_00206_));
 sky130_fd_sc_hd__a22o_1 _06075_ (.A1(net1603),
    .A2(net1048),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net600),
    .X(_00207_));
 sky130_fd_sc_hd__a22o_1 _06076_ (.A1(net1595),
    .A2(net1044),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00208_));
 sky130_fd_sc_hd__a22o_1 _06077_ (.A1(net1587),
    .A2(net1049),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net600),
    .X(_00209_));
 sky130_fd_sc_hd__a22o_1 _06078_ (.A1(net1579),
    .A2(net1044),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00210_));
 sky130_fd_sc_hd__a22o_1 _06079_ (.A1(net1564),
    .A2(net1049),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net600),
    .X(_00212_));
 sky130_fd_sc_hd__a22o_1 _06080_ (.A1(net1556),
    .A2(net1048),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net599),
    .X(_00213_));
 sky130_fd_sc_hd__a22o_1 _06081_ (.A1(net1555),
    .A2(net1048),
    .B1(\u_glbl_reg.reg_12[11] ),
    .B2(net598),
    .X(_00214_));
 sky130_fd_sc_hd__a22o_1 _06082_ (.A1(net1542),
    .A2(net1048),
    .B1(\u_glbl_reg.reg_12[12] ),
    .B2(net598),
    .X(_00215_));
 sky130_fd_sc_hd__xnor2_1 _06083_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[0] ),
    .B(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .Y(_01651_));
 sky130_fd_sc_hd__a21oi_1 _06084_ (.A1(_00244_),
    .A2(_01651_),
    .B1(\u_glbl_reg.u_usbclk.high_count[0] ),
    .Y(_00237_));
 sky130_fd_sc_hd__nand2_1 _06085_ (.A(\u_glbl_reg.u_usbclk.high_count[0] ),
    .B(\u_glbl_reg.u_usbclk.high_count[1] ),
    .Y(_01652_));
 sky130_fd_sc_hd__a21oi_1 _06086_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[0] ),
    .A2(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .B1(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .Y(_01653_));
 sky130_fd_sc_hd__and3_1 _06087_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[0] ),
    .B(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .C(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .X(_01654_));
 sky130_fd_sc_hd__o21a_1 _06088_ (.A1(_01653_),
    .A2(_01654_),
    .B1(_00244_),
    .X(_01655_));
 sky130_fd_sc_hd__a21oi_1 _06089_ (.A1(_01148_),
    .A2(_01652_),
    .B1(_01655_),
    .Y(_00238_));
 sky130_fd_sc_hd__nand2_1 _06090_ (.A(\u_glbl_reg.u_usbclk.high_count[2] ),
    .B(_01148_),
    .Y(_01656_));
 sky130_fd_sc_hd__and3_1 _06091_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .B(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .C(\u_glbl_reg.cfg_usb_clk_ctrl[3] ),
    .X(_01657_));
 sky130_fd_sc_hd__and2_1 _06092_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[0] ),
    .B(_01657_),
    .X(_01658_));
 sky130_fd_sc_hd__nor2_1 _06093_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[3] ),
    .B(_01654_),
    .Y(_01659_));
 sky130_fd_sc_hd__o21a_1 _06094_ (.A1(_01658_),
    .A2(_01659_),
    .B1(_00244_),
    .X(_01660_));
 sky130_fd_sc_hd__a21oi_1 _06095_ (.A1(_01149_),
    .A2(_01656_),
    .B1(_01660_),
    .Y(_00239_));
 sky130_fd_sc_hd__nand2_1 _06096_ (.A(\u_glbl_reg.u_usbclk.high_count[3] ),
    .B(_01149_),
    .Y(_01661_));
 sky130_fd_sc_hd__nor2_1 _06097_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[4] ),
    .B(_01658_),
    .Y(_01662_));
 sky130_fd_sc_hd__and3_1 _06098_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[4] ),
    .B(_00244_),
    .C(_01658_),
    .X(_01663_));
 sky130_fd_sc_hd__a221oi_1 _06099_ (.A1(_01150_),
    .A2(_01661_),
    .B1(_01662_),
    .B2(_00244_),
    .C1(_01663_),
    .Y(_00240_));
 sky130_fd_sc_hd__a21o_1 _06100_ (.A1(\u_glbl_reg.u_usbclk.high_count[4] ),
    .A2(_01150_),
    .B1(_01663_),
    .X(_00241_));
 sky130_fd_sc_hd__a21oi_1 _06101_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .A2(_01155_),
    .B1(\u_glbl_reg.u_usbclk.low_count[0] ),
    .Y(_00245_));
 sky130_fd_sc_hd__and2_1 _06102_ (.A(\u_glbl_reg.u_usbclk.low_count[1] ),
    .B(\u_glbl_reg.u_usbclk.low_count[0] ),
    .X(_01664_));
 sky130_fd_sc_hd__xor2_1 _06103_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .B(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .X(_01665_));
 sky130_fd_sc_hd__o22a_1 _06104_ (.A1(_01151_),
    .A2(_01664_),
    .B1(_01665_),
    .B2(_01156_),
    .X(_00246_));
 sky130_fd_sc_hd__o21ai_1 _06105_ (.A1(\u_glbl_reg.u_usbclk.low_count[1] ),
    .A2(\u_glbl_reg.u_usbclk.low_count[0] ),
    .B1(\u_glbl_reg.u_usbclk.low_count[2] ),
    .Y(_01666_));
 sky130_fd_sc_hd__a21oi_1 _06106_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .A2(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .B1(\u_glbl_reg.cfg_usb_clk_ctrl[3] ),
    .Y(_01667_));
 sky130_fd_sc_hd__nor2_1 _06107_ (.A(_01657_),
    .B(_01667_),
    .Y(_01668_));
 sky130_fd_sc_hd__o2bb2a_1 _06108_ (.A1_N(_01152_),
    .A2_N(_01666_),
    .B1(_01668_),
    .B2(_01156_),
    .X(_00247_));
 sky130_fd_sc_hd__and2_1 _06109_ (.A(\u_glbl_reg.u_usbclk.low_count[3] ),
    .B(_01152_),
    .X(_01669_));
 sky130_fd_sc_hd__xor2_1 _06110_ (.A(\u_glbl_reg.cfg_usb_clk_ctrl[4] ),
    .B(_01657_),
    .X(_01670_));
 sky130_fd_sc_hd__o22a_1 _06111_ (.A1(_01154_),
    .A2(_01669_),
    .B1(_01670_),
    .B2(_01156_),
    .X(_00248_));
 sky130_fd_sc_hd__and2_1 _06112_ (.A(\u_glbl_reg.u_usbclk.low_count[4] ),
    .B(_01153_),
    .X(_01671_));
 sky130_fd_sc_hd__a31o_1 _06113_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[4] ),
    .A2(_01155_),
    .A3(_01657_),
    .B1(_01671_),
    .X(_00249_));
 sky130_fd_sc_hd__mux2_1 _06114_ (.A0(clknet_1_0__leaf_user_clock1),
    .A1(clknet_1_1__leaf_user_clock2),
    .S(\u_glbl_reg.cfg_rtc_clk_ctrl[6] ),
    .X(_01672_));
 sky130_fd_sc_hd__mux2_1 _06115_ (.A0(_01672_),
    .A1(net1375),
    .S(\u_glbl_reg.cfg_rtc_clk_ctrl[7] ),
    .X(\u_glbl_reg.rtc_ref_clk_int ));
 sky130_fd_sc_hd__mux2_1 _06116_ (.A0(clknet_1_0__leaf_user_clock1),
    .A1(clknet_1_0__leaf_user_clock2),
    .S(\u_glbl_reg.cfg_usb_clk_ctrl[6] ),
    .X(_01673_));
 sky130_fd_sc_hd__mux2_1 _06117_ (.A0(_01673_),
    .A1(net1375),
    .S(\u_glbl_reg.cfg_usb_clk_ctrl[7] ),
    .X(\u_glbl_reg.u_usb_ref_clkbuf.A ));
 sky130_fd_sc_hd__mux4_2 _06118_ (.A0(clknet_1_0__leaf_user_clock1),
    .A1(clknet_1_0__leaf_user_clock2),
    .A2(net1375),
    .A3(net45),
    .S0(\u_glbl_reg.cfg_mon_sel[0] ),
    .S1(\u_glbl_reg.cfg_mon_sel[1] ),
    .X(_01674_));
 sky130_fd_sc_hd__mux4_2 _06119_ (.A0(clknet_leaf_118_mclk),
    .A1(net2),
    .A2(net504),
    .A3(net454),
    .S0(\u_glbl_reg.cfg_mon_sel[0] ),
    .S1(\u_glbl_reg.cfg_mon_sel[1] ),
    .X(_01675_));
 sky130_fd_sc_hd__inv_2 _06120__1 (.A(_01675_),
    .Y(net1691));
 sky130_fd_sc_hd__a21oi_2 _06121_ (.A1(\u_glbl_reg.cfg_mon_sel[2] ),
    .A2(net1691),
    .B1(\u_glbl_reg.cfg_mon_sel[3] ),
    .Y(_01677_));
 sky130_fd_sc_hd__o21a_2 _06122_ (.A1(\u_glbl_reg.cfg_mon_sel[2] ),
    .A2(_01674_),
    .B1(_01677_),
    .X(\u_glbl_reg.dbg_clk_ref ));
 sky130_fd_sc_hd__or2_1 _06123_ (.A(net1293),
    .B(net1202),
    .X(_00091_));
 sky130_fd_sc_hd__or2_1 _06124_ (.A(net1572),
    .B(net1201),
    .X(_00102_));
 sky130_fd_sc_hd__and2b_1 _06125_ (.A_N(net1201),
    .B(net1488),
    .X(_00113_));
 sky130_fd_sc_hd__and2b_1 _06126_ (.A_N(net1202),
    .B(net1466),
    .X(_00116_));
 sky130_fd_sc_hd__and2b_1 _06127_ (.A_N(net1202),
    .B(net1457),
    .X(_00117_));
 sky130_fd_sc_hd__and2b_1 _06128_ (.A_N(net1201),
    .B(net1448),
    .X(_00118_));
 sky130_fd_sc_hd__and2b_1 _06129_ (.A_N(net1201),
    .B(net1441),
    .X(_00119_));
 sky130_fd_sc_hd__and2b_1 _06130_ (.A_N(net1201),
    .B(net1433),
    .X(_00120_));
 sky130_fd_sc_hd__a22o_1 _06131_ (.A1(\u_gpio.u_bit[0].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[0] ),
    .X(_01678_));
 sky130_fd_sc_hd__a221o_1 _06132_ (.A1(\u_gpio.cfg_gpio_out_type[0] ),
    .A2(net704),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[0] ),
    .C1(_01678_),
    .X(_01679_));
 sky130_fd_sc_hd__a221o_1 _06133_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[0] ),
    .A2(net670),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[0] ),
    .C1(_01679_),
    .X(_01680_));
 sky130_fd_sc_hd__a221o_1 _06134_ (.A1(net1814),
    .A2(net717),
    .B1(net667),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[0] ),
    .C1(_01680_),
    .X(\u_gpio.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__a22o_1 _06135_ (.A1(\u_gpio.cfg_gpio_out_data[1] ),
    .A2(net1138),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[1] ),
    .X(_01681_));
 sky130_fd_sc_hd__a221o_1 _06136_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.data_out ),
    .A2(net715),
    .B1(net692),
    .B2(net1844),
    .C1(_01681_),
    .X(_01682_));
 sky130_fd_sc_hd__a22o_1 _06137_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[1] ),
    .A2(net668),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[1] ),
    .X(_01683_));
 sky130_fd_sc_hd__a221o_1 _06138_ (.A1(\u_gpio.cfg_gpio_out_type[1] ),
    .A2(net704),
    .B1(net664),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[1] ),
    .C1(_01683_),
    .X(_01684_));
 sky130_fd_sc_hd__or2_1 _06139_ (.A(net1845),
    .B(_01684_),
    .X(\u_gpio.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__a22o_1 _06140_ (.A1(\u_gpio.cfg_gpio_out_type[2] ),
    .A2(net704),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[2] ),
    .X(_01685_));
 sky130_fd_sc_hd__a221o_1 _06141_ (.A1(\u_gpio.u_bit[2].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[2] ),
    .C1(_01685_),
    .X(_01686_));
 sky130_fd_sc_hd__a221o_1 _06142_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[2] ),
    .A2(net670),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[2] ),
    .C1(_01686_),
    .X(_01687_));
 sky130_fd_sc_hd__a221o_1 _06143_ (.A1(net1818),
    .A2(net717),
    .B1(net667),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[2] ),
    .C1(_01687_),
    .X(\u_gpio.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__a22o_1 _06144_ (.A1(\u_gpio.cfg_gpio_out_type[3] ),
    .A2(net704),
    .B1(net1141),
    .B2(\u_gpio.cfg_gpio_out_data[3] ),
    .X(_01688_));
 sky130_fd_sc_hd__a221o_1 _06145_ (.A1(net1831),
    .A2(net692),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[3] ),
    .C1(_01688_),
    .X(_01689_));
 sky130_fd_sc_hd__a22o_1 _06146_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.data_out ),
    .A2(net716),
    .B1(net668),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[3] ),
    .X(_01690_));
 sky130_fd_sc_hd__a221o_1 _06147_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[3] ),
    .A2(net664),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[3] ),
    .C1(_01690_),
    .X(_01691_));
 sky130_fd_sc_hd__or2_1 _06148_ (.A(net1832),
    .B(_01691_),
    .X(\u_gpio.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__a22o_1 _06149_ (.A1(\u_gpio.u_bit[4].u_dglitch.gpio_reg ),
    .A2(net692),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[4] ),
    .X(_01692_));
 sky130_fd_sc_hd__a221o_1 _06150_ (.A1(\u_gpio.cfg_gpio_out_type[4] ),
    .A2(net704),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[4] ),
    .C1(_01692_),
    .X(_01693_));
 sky130_fd_sc_hd__a221o_1 _06151_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[4] ),
    .A2(_01538_),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[4] ),
    .C1(_01693_),
    .X(_01694_));
 sky130_fd_sc_hd__a221o_1 _06152_ (.A1(net1820),
    .A2(net716),
    .B1(net664),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[4] ),
    .C1(_01694_),
    .X(\u_gpio.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__a22o_1 _06153_ (.A1(net1828),
    .A2(net717),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[5] ),
    .X(_01695_));
 sky130_fd_sc_hd__a22o_1 _06154_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[5] ),
    .A2(net668),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[5] ),
    .X(_01696_));
 sky130_fd_sc_hd__a221o_1 _06155_ (.A1(\u_gpio.cfg_gpio_out_type[5] ),
    .A2(net704),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[5] ),
    .C1(_01696_),
    .X(_01697_));
 sky130_fd_sc_hd__a211o_1 _06156_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[5] ),
    .A2(net667),
    .B1(net1829),
    .C1(_01697_),
    .X(\u_gpio.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__and3_1 _06157_ (.A(\u_gpio.cfg_gpio_negedge_int_sel[6] ),
    .B(net1242),
    .C(net1153),
    .X(_01698_));
 sky130_fd_sc_hd__a22o_1 _06158_ (.A1(net1847),
    .A2(net717),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[6] ),
    .X(_01699_));
 sky130_fd_sc_hd__a221o_1 _06159_ (.A1(\u_gpio.cfg_gpio_out_type[6] ),
    .A2(net704),
    .B1(net670),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[6] ),
    .C1(_01698_),
    .X(_01700_));
 sky130_fd_sc_hd__a22o_1 _06160_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[6] ),
    .A2(net664),
    .B1(net1133),
    .B2(\u_gpio.cfg_gpio_dir_sel[6] ),
    .X(_01701_));
 sky130_fd_sc_hd__or3_1 _06161_ (.A(net1848),
    .B(_01700_),
    .C(_01701_),
    .X(\u_gpio.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__a22o_1 _06162_ (.A1(net1836),
    .A2(net715),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[7] ),
    .X(_01702_));
 sky130_fd_sc_hd__a22o_1 _06163_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[7] ),
    .A2(net668),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[7] ),
    .X(_01703_));
 sky130_fd_sc_hd__a221o_1 _06164_ (.A1(\u_gpio.cfg_gpio_out_type[7] ),
    .A2(net704),
    .B1(_01539_),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[7] ),
    .C1(_01703_),
    .X(_01704_));
 sky130_fd_sc_hd__a211o_1 _06165_ (.A1(\u_gpio.cfg_gpio_dir_sel[7] ),
    .A2(net1133),
    .B1(net1837),
    .C1(_01704_),
    .X(\u_gpio.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__a22o_1 _06166_ (.A1(\u_gpio.cfg_gpio_out_type[8] ),
    .A2(net703),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[8] ),
    .X(_01705_));
 sky130_fd_sc_hd__a221o_1 _06167_ (.A1(\u_gpio.u_bit[8].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[8] ),
    .C1(_01705_),
    .X(_01706_));
 sky130_fd_sc_hd__a221o_1 _06168_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[8] ),
    .A2(net667),
    .B1(net1137),
    .B2(\u_gpio.cfg_gpio_out_data[8] ),
    .C1(_01706_),
    .X(_01707_));
 sky130_fd_sc_hd__a221o_1 _06169_ (.A1(net1868),
    .A2(net717),
    .B1(net670),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[8] ),
    .C1(_01707_),
    .X(\u_gpio.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__a22o_1 _06170_ (.A1(\u_gpio.cfg_gpio_dir_sel[9] ),
    .A2(net1132),
    .B1(net663),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[9] ),
    .X(_01708_));
 sky130_fd_sc_hd__a221o_1 _06171_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.data_out ),
    .A2(net716),
    .B1(net691),
    .B2(net1850),
    .C1(_01708_),
    .X(_01709_));
 sky130_fd_sc_hd__a22o_1 _06172_ (.A1(\u_gpio.cfg_gpio_out_type[9] ),
    .A2(net702),
    .B1(net664),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[9] ),
    .X(_01710_));
 sky130_fd_sc_hd__a221o_1 _06173_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[9] ),
    .A2(net668),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[9] ),
    .C1(_01710_),
    .X(_01711_));
 sky130_fd_sc_hd__or2_2 _06174_ (.A(net1851),
    .B(_01711_),
    .X(\u_gpio.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__a22o_1 _06175_ (.A1(\u_gpio.cfg_gpio_out_type[10] ),
    .A2(net702),
    .B1(net664),
    .B2(\u_gpio.u_reg.cfg_gpio_int_mask[10] ),
    .X(_01712_));
 sky130_fd_sc_hd__a221o_1 _06176_ (.A1(\u_gpio.cfg_gpio_out_data[10] ),
    .A2(net1136),
    .B1(net663),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[10] ),
    .C1(_01712_),
    .X(_01713_));
 sky130_fd_sc_hd__a22o_1 _06177_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.data_out ),
    .A2(net716),
    .B1(net691),
    .B2(net1998),
    .X(_01714_));
 sky130_fd_sc_hd__a221o_1 _06178_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[10] ),
    .A2(net668),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[10] ),
    .C1(net1999),
    .X(_01715_));
 sky130_fd_sc_hd__or2_1 _06179_ (.A(_01713_),
    .B(_01715_),
    .X(\u_gpio.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__a22o_1 _06180_ (.A1(\u_gpio.u_bit[11].u_dglitch.gpio_reg ),
    .A2(net692),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[11] ),
    .X(_01716_));
 sky130_fd_sc_hd__a221o_1 _06181_ (.A1(\u_gpio.cfg_gpio_out_type[11] ),
    .A2(net702),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[11] ),
    .C1(_01716_),
    .X(_01717_));
 sky130_fd_sc_hd__a221o_1 _06182_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[11] ),
    .A2(net664),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[11] ),
    .C1(_01717_),
    .X(_01718_));
 sky130_fd_sc_hd__a221o_1 _06183_ (.A1(net1878),
    .A2(net716),
    .B1(net668),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[11] ),
    .C1(_01718_),
    .X(\u_gpio.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__a22o_1 _06184_ (.A1(\u_gpio.cfg_gpio_out_type[12] ),
    .A2(net703),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[12] ),
    .X(_01719_));
 sky130_fd_sc_hd__a221o_1 _06185_ (.A1(\u_gpio.u_bit[12].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[12] ),
    .C1(_01719_),
    .X(_01720_));
 sky130_fd_sc_hd__a221o_1 _06186_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[12] ),
    .A2(net664),
    .B1(net1137),
    .B2(\u_gpio.cfg_gpio_out_data[12] ),
    .C1(_01720_),
    .X(_01721_));
 sky130_fd_sc_hd__a221o_1 _06187_ (.A1(net1899),
    .A2(net716),
    .B1(net668),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[12] ),
    .C1(_01721_),
    .X(\u_gpio.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__a22o_1 _06188_ (.A1(\u_gpio.cfg_gpio_out_type[13] ),
    .A2(net703),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[13] ),
    .X(_01722_));
 sky130_fd_sc_hd__a221o_1 _06189_ (.A1(\u_gpio.u_bit[13].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[13] ),
    .C1(_01722_),
    .X(_01723_));
 sky130_fd_sc_hd__a221o_1 _06190_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[13] ),
    .A2(net664),
    .B1(net1137),
    .B2(\u_gpio.cfg_gpio_out_data[13] ),
    .C1(_01723_),
    .X(_01724_));
 sky130_fd_sc_hd__a221o_1 _06191_ (.A1(net1895),
    .A2(net716),
    .B1(net668),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[13] ),
    .C1(_01724_),
    .X(\u_gpio.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__a22o_1 _06192_ (.A1(\u_gpio.cfg_gpio_out_type[14] ),
    .A2(net703),
    .B1(net1137),
    .B2(\u_gpio.cfg_gpio_out_data[14] ),
    .X(_01725_));
 sky130_fd_sc_hd__a221o_1 _06193_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[14] ),
    .A2(net667),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[14] ),
    .C1(_01725_),
    .X(_01726_));
 sky130_fd_sc_hd__a22o_1 _06194_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.data_out ),
    .A2(net717),
    .B1(net693),
    .B2(net1933),
    .X(_01727_));
 sky130_fd_sc_hd__a221o_1 _06195_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[14] ),
    .A2(net670),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[14] ),
    .C1(net1934),
    .X(_01728_));
 sky130_fd_sc_hd__or2_1 _06196_ (.A(_01726_),
    .B(net1935),
    .X(\u_gpio.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__a22o_1 _06197_ (.A1(\u_gpio.u_bit[15].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[15] ),
    .X(_01729_));
 sky130_fd_sc_hd__a221o_1 _06198_ (.A1(\u_gpio.cfg_gpio_out_type[15] ),
    .A2(net703),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[15] ),
    .C1(_01729_),
    .X(_01730_));
 sky130_fd_sc_hd__a221o_1 _06199_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[15] ),
    .A2(net667),
    .B1(net1137),
    .B2(\u_gpio.cfg_gpio_out_data[15] ),
    .C1(_01730_),
    .X(_01731_));
 sky130_fd_sc_hd__a221o_1 _06200_ (.A1(net1953),
    .A2(net717),
    .B1(net670),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[15] ),
    .C1(_01731_),
    .X(\u_gpio.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__a22o_1 _06201_ (.A1(\u_gpio.u_bit[16].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net662),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[16] ),
    .X(_01732_));
 sky130_fd_sc_hd__a221o_1 _06202_ (.A1(\u_gpio.cfg_gpio_out_type[16] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[16] ),
    .C1(_01732_),
    .X(_01733_));
 sky130_fd_sc_hd__a221o_1 _06203_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[16] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[16] ),
    .C1(_01733_),
    .X(_01734_));
 sky130_fd_sc_hd__a221o_1 _06204_ (.A1(net1861),
    .A2(net717),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[16] ),
    .C1(_01734_),
    .X(\u_gpio.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__a22o_1 _06205_ (.A1(\u_gpio.u_bit[17].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net662),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[17] ),
    .X(_01735_));
 sky130_fd_sc_hd__a221o_1 _06206_ (.A1(\u_gpio.cfg_gpio_out_type[17] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[17] ),
    .C1(_01735_),
    .X(_01736_));
 sky130_fd_sc_hd__a221o_1 _06207_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[17] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[17] ),
    .C1(_01736_),
    .X(_01737_));
 sky130_fd_sc_hd__a221o_1 _06208_ (.A1(net1957),
    .A2(net717),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[17] ),
    .C1(_01737_),
    .X(\u_gpio.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__a22o_1 _06209_ (.A1(\u_gpio.cfg_gpio_out_type[18] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[18] ),
    .X(_01738_));
 sky130_fd_sc_hd__a221o_1 _06210_ (.A1(\u_gpio.u_bit[18].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[18] ),
    .C1(_01738_),
    .X(_01739_));
 sky130_fd_sc_hd__a221o_1 _06211_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[18] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[18] ),
    .C1(_01739_),
    .X(_01740_));
 sky130_fd_sc_hd__a221o_1 _06212_ (.A1(net1951),
    .A2(net718),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[18] ),
    .C1(_01740_),
    .X(\u_gpio.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__a22o_1 _06213_ (.A1(\u_gpio.u_bit[19].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[19] ),
    .X(_01741_));
 sky130_fd_sc_hd__a221o_1 _06214_ (.A1(\u_gpio.cfg_gpio_out_type[19] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[19] ),
    .C1(_01741_),
    .X(_01742_));
 sky130_fd_sc_hd__a221o_1 _06215_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[19] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[19] ),
    .C1(_01742_),
    .X(_01743_));
 sky130_fd_sc_hd__a221o_1 _06216_ (.A1(net1946),
    .A2(net718),
    .B1(net670),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[19] ),
    .C1(_01743_),
    .X(\u_gpio.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__a22o_1 _06217_ (.A1(\u_gpio.cfg_gpio_out_type[20] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[20] ),
    .X(_01744_));
 sky130_fd_sc_hd__a221o_1 _06218_ (.A1(\u_gpio.u_bit[20].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[20] ),
    .C1(_01744_),
    .X(_01745_));
 sky130_fd_sc_hd__a221o_1 _06219_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[20] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[20] ),
    .C1(_01745_),
    .X(_01746_));
 sky130_fd_sc_hd__a221o_1 _06220_ (.A1(net1941),
    .A2(net718),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[20] ),
    .C1(_01746_),
    .X(\u_gpio.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__a22o_1 _06221_ (.A1(\u_gpio.u_bit[21].u_dglitch.gpio_reg ),
    .A2(net697),
    .B1(net662),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[21] ),
    .X(_01747_));
 sky130_fd_sc_hd__a221o_1 _06222_ (.A1(\u_gpio.cfg_gpio_out_type[21] ),
    .A2(net707),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[21] ),
    .C1(_01747_),
    .X(_01748_));
 sky130_fd_sc_hd__a221o_1 _06223_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[21] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[21] ),
    .C1(_01748_),
    .X(_01749_));
 sky130_fd_sc_hd__a221o_1 _06224_ (.A1(net1955),
    .A2(net718),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[21] ),
    .C1(_01749_),
    .X(\u_gpio.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__a22o_1 _06225_ (.A1(\u_gpio.cfg_gpio_out_type[22] ),
    .A2(net703),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[22] ),
    .X(_01750_));
 sky130_fd_sc_hd__a221o_1 _06226_ (.A1(\u_gpio.u_bit[22].u_dglitch.gpio_reg ),
    .A2(net693),
    .B1(net1134),
    .B2(\u_gpio.cfg_gpio_dir_sel[22] ),
    .C1(_01750_),
    .X(_01751_));
 sky130_fd_sc_hd__a221o_1 _06227_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[22] ),
    .A2(net666),
    .B1(net1139),
    .B2(\u_gpio.cfg_gpio_out_data[22] ),
    .C1(_01751_),
    .X(_01752_));
 sky130_fd_sc_hd__a221o_1 _06228_ (.A1(net1962),
    .A2(net717),
    .B1(net671),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[22] ),
    .C1(_01752_),
    .X(\u_gpio.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__a22o_1 _06229_ (.A1(\u_gpio.cfg_gpio_out_type[23] ),
    .A2(net707),
    .B1(net670),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[23] ),
    .X(_01753_));
 sky130_fd_sc_hd__a22o_1 _06230_ (.A1(\u_gpio.cfg_gpio_dir_sel[23] ),
    .A2(net1134),
    .B1(net661),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[23] ),
    .X(_01754_));
 sky130_fd_sc_hd__a221o_1 _06231_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[23] ),
    .A2(net666),
    .B1(net1140),
    .B2(\u_gpio.cfg_gpio_out_data[23] ),
    .C1(_01753_),
    .X(_01755_));
 sky130_fd_sc_hd__a211o_1 _06232_ (.A1(net1943),
    .A2(net718),
    .B1(_01754_),
    .C1(_01755_),
    .X(\u_gpio.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__a22o_1 _06233_ (.A1(\u_gpio.u_bit[24].u_dglitch.gpio_reg ),
    .A2(net691),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[24] ),
    .X(_01756_));
 sky130_fd_sc_hd__a221o_1 _06234_ (.A1(\u_gpio.cfg_gpio_out_type[24] ),
    .A2(net702),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[24] ),
    .C1(_01756_),
    .X(_01757_));
 sky130_fd_sc_hd__a221o_1 _06235_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[24] ),
    .A2(net665),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[24] ),
    .C1(_01757_),
    .X(_01758_));
 sky130_fd_sc_hd__a221o_1 _06236_ (.A1(net1949),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[24] ),
    .C1(_01758_),
    .X(\u_gpio.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__a22o_1 _06237_ (.A1(\u_gpio.cfg_gpio_out_type[25] ),
    .A2(net702),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[25] ),
    .X(_01759_));
 sky130_fd_sc_hd__a221o_1 _06238_ (.A1(net1922),
    .A2(net691),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[25] ),
    .C1(_01759_),
    .X(_01760_));
 sky130_fd_sc_hd__a221o_1 _06239_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[25] ),
    .A2(net665),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[25] ),
    .C1(net1923),
    .X(_01761_));
 sky130_fd_sc_hd__a221o_1 _06240_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.data_out ),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[25] ),
    .C1(net1924),
    .X(\u_gpio.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__a22o_1 _06241_ (.A1(\u_gpio.cfg_gpio_out_type[26] ),
    .A2(net702),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[26] ),
    .X(_01762_));
 sky130_fd_sc_hd__a221o_1 _06242_ (.A1(\u_gpio.u_bit[26].u_dglitch.gpio_reg ),
    .A2(net691),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[26] ),
    .C1(_01762_),
    .X(_01763_));
 sky130_fd_sc_hd__a221o_1 _06243_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[26] ),
    .A2(net665),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[26] ),
    .C1(_01763_),
    .X(_01764_));
 sky130_fd_sc_hd__a221o_1 _06244_ (.A1(net1937),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[26] ),
    .C1(_01764_),
    .X(\u_gpio.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__a22o_1 _06245_ (.A1(\u_gpio.cfg_gpio_out_type[27] ),
    .A2(net703),
    .B1(net660),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[27] ),
    .X(_01765_));
 sky130_fd_sc_hd__a221o_1 _06246_ (.A1(\u_gpio.u_bit[27].u_dglitch.gpio_reg ),
    .A2(net691),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[27] ),
    .C1(_01765_),
    .X(_01766_));
 sky130_fd_sc_hd__a221o_1 _06247_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[27] ),
    .A2(net665),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[27] ),
    .C1(_01766_),
    .X(_01767_));
 sky130_fd_sc_hd__a221o_1 _06248_ (.A1(net1910),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[27] ),
    .C1(_01767_),
    .X(\u_gpio.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__a22o_1 _06249_ (.A1(\u_gpio.cfg_gpio_out_type[28] ),
    .A2(net703),
    .B1(net1138),
    .B2(\u_gpio.cfg_gpio_out_data[28] ),
    .X(_01768_));
 sky130_fd_sc_hd__a221o_1 _06250_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[28] ),
    .A2(net665),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[28] ),
    .C1(_01768_),
    .X(_01769_));
 sky130_fd_sc_hd__a22o_1 _06251_ (.A1(net1839),
    .A2(net715),
    .B1(net691),
    .B2(\u_gpio.u_bit[28].u_dglitch.gpio_reg ),
    .X(_01770_));
 sky130_fd_sc_hd__a221o_1 _06252_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[28] ),
    .A2(net669),
    .B1(net1132),
    .B2(\u_gpio.cfg_gpio_dir_sel[28] ),
    .C1(net1840),
    .X(_01771_));
 sky130_fd_sc_hd__or2_1 _06253_ (.A(_01769_),
    .B(net1841),
    .X(\u_gpio.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__a22o_1 _06254_ (.A1(\u_gpio.cfg_gpio_out_type[29] ),
    .A2(net703),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[29] ),
    .X(_01772_));
 sky130_fd_sc_hd__a221o_1 _06255_ (.A1(\u_gpio.u_bit[29].u_dglitch.gpio_reg ),
    .A2(net691),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[29] ),
    .C1(_01772_),
    .X(_01773_));
 sky130_fd_sc_hd__a221o_1 _06256_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[29] ),
    .A2(net665),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[29] ),
    .C1(_01773_),
    .X(_01774_));
 sky130_fd_sc_hd__a221o_1 _06257_ (.A1(net1944),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[29] ),
    .C1(_01774_),
    .X(\u_gpio.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__a22o_1 _06258_ (.A1(\u_gpio.cfg_gpio_out_type[30] ),
    .A2(net702),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[30] ),
    .X(_01775_));
 sky130_fd_sc_hd__a221o_1 _06259_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[30] ),
    .A2(net665),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[30] ),
    .C1(_01775_),
    .X(_01776_));
 sky130_fd_sc_hd__a22o_1 _06260_ (.A1(\u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.data_out ),
    .A2(net715),
    .B1(net691),
    .B2(net1978),
    .X(_01777_));
 sky130_fd_sc_hd__a221o_1 _06261_ (.A1(\u_gpio.cfg_gpio_posedge_int_sel[30] ),
    .A2(net669),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[30] ),
    .C1(net1979),
    .X(_01778_));
 sky130_fd_sc_hd__or2_1 _06262_ (.A(_01776_),
    .B(net1980),
    .X(\u_gpio.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__a22o_1 _06263_ (.A1(\u_gpio.cfg_gpio_out_type[31] ),
    .A2(net702),
    .B1(net659),
    .B2(\u_gpio.cfg_gpio_negedge_int_sel[31] ),
    .X(_01779_));
 sky130_fd_sc_hd__a221o_1 _06264_ (.A1(\u_gpio.u_bit[31].u_dglitch.gpio_reg ),
    .A2(net691),
    .B1(net1131),
    .B2(\u_gpio.cfg_gpio_dir_sel[31] ),
    .C1(_01779_),
    .X(_01780_));
 sky130_fd_sc_hd__a221o_1 _06265_ (.A1(\u_gpio.u_reg.cfg_gpio_int_mask[31] ),
    .A2(net665),
    .B1(net1136),
    .B2(\u_gpio.cfg_gpio_out_data[31] ),
    .C1(_01780_),
    .X(_01781_));
 sky130_fd_sc_hd__a221o_1 _06266_ (.A1(net1920),
    .A2(net715),
    .B1(net669),
    .B2(\u_gpio.cfg_gpio_posedge_int_sel[31] ),
    .C1(_01781_),
    .X(\u_gpio.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__nor2_2 _06267_ (.A(net1225),
    .B(_01145_),
    .Y(_01782_));
 sky130_fd_sc_hd__a22o_1 _06268_ (.A1(\u_glbl_reg.reg_3[0] ),
    .A2(net621),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[0] ),
    .X(_01783_));
 sky130_fd_sc_hd__a221o_1 _06269_ (.A1(\u_glbl_reg.reg_20[0] ),
    .A2(net638),
    .B1(net608),
    .B2(\u_glbl_reg.cfg_ref_pll_div[0] ),
    .C1(_01783_),
    .X(_01784_));
 sky130_fd_sc_hd__a22o_1 _06270_ (.A1(net1254),
    .A2(net711),
    .B1(net1161),
    .B2(_01118_),
    .X(_01785_));
 sky130_fd_sc_hd__and3_4 _06271_ (.A(net1254),
    .B(net1247),
    .C(net1214),
    .X(_01786_));
 sky130_fd_sc_hd__a221o_1 _06272_ (.A1(\u_glbl_reg.reg_18[0] ),
    .A2(net646),
    .B1(net561),
    .B2(net2317),
    .C1(_01786_),
    .X(_01787_));
 sky130_fd_sc_hd__and3_1 _06273_ (.A(net1254),
    .B(net1179),
    .C(net1153),
    .X(_01788_));
 sky130_fd_sc_hd__nand2_8 _06274_ (.A(net1179),
    .B(_01118_),
    .Y(_01789_));
 sky130_fd_sc_hd__nand2_2 _06275_ (.A(\u_glbl_reg.u_random.n1_plus_n0[15] ),
    .B(\u_glbl_reg.u_random.n0[0] ),
    .Y(_01790_));
 sky130_fd_sc_hd__or2_1 _06276_ (.A(\u_glbl_reg.u_random.n1_plus_n0[15] ),
    .B(\u_glbl_reg.u_random.n0[0] ),
    .X(_01791_));
 sky130_fd_sc_hd__a32o_4 _06277_ (.A1(net594),
    .A2(_01790_),
    .A3(_01791_),
    .B1(net606),
    .B2(net199),
    .X(_01792_));
 sky130_fd_sc_hd__nor2_4 _06278_ (.A(_01115_),
    .B(_01145_),
    .Y(_01793_));
 sky130_fd_sc_hd__a221o_1 _06279_ (.A1(net465),
    .A2(net682),
    .B1(net590),
    .B2(net159),
    .C1(_01792_),
    .X(_01794_));
 sky130_fd_sc_hd__a22o_1 _06280_ (.A1(\u_glbl_reg.reg_17[0] ),
    .A2(net649),
    .B1(net624),
    .B2(\u_glbl_reg.reg_23[0] ),
    .X(_01795_));
 sky130_fd_sc_hd__a221o_1 _06281_ (.A1(\u_glbl_reg.reg_22[0] ),
    .A2(net628),
    .B1(net617),
    .B2(\u_glbl_reg.cfg_multi_func_sel[0] ),
    .C1(_01795_),
    .X(_01796_));
 sky130_fd_sc_hd__and2_1 _06282_ (.A(\u_glbl_reg.reg_21[0] ),
    .B(net634),
    .X(_01797_));
 sky130_fd_sc_hd__a221o_1 _06283_ (.A1(\u_glbl_reg.reg_15[0] ),
    .A2(net655),
    .B1(net1125),
    .B2(\u_glbl_reg.reg_16[0] ),
    .C1(_01797_),
    .X(_01798_));
 sky130_fd_sc_hd__a22o_1 _06284_ (.A1(\u_glbl_reg.reg_2[0] ),
    .A2(net686),
    .B1(net642),
    .B2(\u_glbl_reg.reg_19[0] ),
    .X(_01799_));
 sky130_fd_sc_hd__a221o_1 _06285_ (.A1(\u_glbl_reg.cfg_rst_ctrl[0] ),
    .A2(net698),
    .B1(net613),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ),
    .C1(_01799_),
    .X(_01800_));
 sky130_fd_sc_hd__or4_1 _06286_ (.A(_01794_),
    .B(_01796_),
    .C(_01798_),
    .D(_01800_),
    .X(_01801_));
 sky130_fd_sc_hd__or3_2 _06287_ (.A(_01784_),
    .B(_01787_),
    .C(_01801_),
    .X(\u_glbl_reg.reg_out[0] ));
 sky130_fd_sc_hd__nand2_1 _06288_ (.A(\u_glbl_reg.u_random.n1_plus_n0[16] ),
    .B(\u_glbl_reg.u_random.n0[1] ),
    .Y(_01802_));
 sky130_fd_sc_hd__nor2_1 _06289_ (.A(\u_glbl_reg.u_random.n1_plus_n0[16] ),
    .B(\u_glbl_reg.u_random.n0[1] ),
    .Y(_01803_));
 sky130_fd_sc_hd__or2_1 _06290_ (.A(\u_glbl_reg.u_random.n1_plus_n0[16] ),
    .B(\u_glbl_reg.u_random.n0[1] ),
    .X(_01804_));
 sky130_fd_sc_hd__a21bo_2 _06291_ (.A1(_01802_),
    .A2(_01804_),
    .B1_N(_01790_),
    .X(_01805_));
 sky130_fd_sc_hd__and3b_1 _06292_ (.A_N(_01790_),
    .B(_01802_),
    .C(_01804_),
    .X(_01806_));
 sky130_fd_sc_hd__inv_2 _06293_ (.A(_01806_),
    .Y(_01807_));
 sky130_fd_sc_hd__a22o_1 _06294_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ),
    .A2(net613),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[1] ),
    .X(_01808_));
 sky130_fd_sc_hd__a22o_1 _06295_ (.A1(\u_glbl_reg.reg_23[1] ),
    .A2(net625),
    .B1(net608),
    .B2(\u_glbl_reg.cfg_ref_pll_div[1] ),
    .X(_01809_));
 sky130_fd_sc_hd__a22o_1 _06296_ (.A1(\u_glbl_reg.reg_17[1] ),
    .A2(net650),
    .B1(net590),
    .B2(net170),
    .X(_01810_));
 sky130_fd_sc_hd__a221o_1 _06297_ (.A1(\u_glbl_reg.reg_18[1] ),
    .A2(net646),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[1] ),
    .C1(_01810_),
    .X(_01811_));
 sky130_fd_sc_hd__a221o_1 _06298_ (.A1(\u_glbl_reg.reg_2[1] ),
    .A2(net686),
    .B1(net654),
    .B2(\u_glbl_reg.reg_15[1] ),
    .C1(_01808_),
    .X(_01812_));
 sky130_fd_sc_hd__a221o_1 _06299_ (.A1(net2062),
    .A2(net1124),
    .B1(net642),
    .B2(\u_glbl_reg.reg_19[1] ),
    .C1(_01809_),
    .X(_01813_));
 sky130_fd_sc_hd__a22o_1 _06300_ (.A1(net476),
    .A2(net683),
    .B1(net621),
    .B2(\u_glbl_reg.reg_3[1] ),
    .X(_01814_));
 sky130_fd_sc_hd__a221o_1 _06301_ (.A1(\u_glbl_reg.cfg_rst_ctrl[1] ),
    .A2(net699),
    .B1(net603),
    .B2(net1099),
    .C1(_01814_),
    .X(_01815_));
 sky130_fd_sc_hd__a32o_1 _06302_ (.A1(net595),
    .A2(_01805_),
    .A3(_01807_),
    .B1(net638),
    .B2(\u_glbl_reg.reg_20[1] ),
    .X(_01816_));
 sky130_fd_sc_hd__a221o_1 _06303_ (.A1(\u_glbl_reg.reg_21[1] ),
    .A2(net634),
    .B1(net619),
    .B2(\u_glbl_reg.cfg_multi_func_sel[1] ),
    .C1(_01816_),
    .X(_01817_));
 sky130_fd_sc_hd__a211o_1 _06304_ (.A1(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ),
    .A2(net561),
    .B1(_01811_),
    .C1(_01815_),
    .X(_01818_));
 sky130_fd_sc_hd__or4_4 _06305_ (.A(_01812_),
    .B(_01813_),
    .C(_01817_),
    .D(_01818_),
    .X(\u_glbl_reg.reg_out[1] ));
 sky130_fd_sc_hd__a22o_1 _06306_ (.A1(\u_glbl_reg.reg_17[2] ),
    .A2(net649),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[2] ),
    .X(_01819_));
 sky130_fd_sc_hd__a221o_1 _06307_ (.A1(\u_glbl_reg.reg_18[2] ),
    .A2(net645),
    .B1(net617),
    .B2(\u_glbl_reg.cfg_multi_func_sel[2] ),
    .C1(_01819_),
    .X(_01820_));
 sky130_fd_sc_hd__a22o_1 _06308_ (.A1(\u_glbl_reg.cfg_rst_ctrl[2] ),
    .A2(net698),
    .B1(net634),
    .B2(\u_glbl_reg.reg_21[2] ),
    .X(_01821_));
 sky130_fd_sc_hd__a221o_1 _06309_ (.A1(\u_glbl_reg.reg_20[2] ),
    .A2(net637),
    .B1(net590),
    .B2(net181),
    .C1(_01821_),
    .X(_01822_));
 sky130_fd_sc_hd__a22o_1 _06310_ (.A1(\u_glbl_reg.reg_2[2] ),
    .A2(net686),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[2] ),
    .X(_01823_));
 sky130_fd_sc_hd__a21o_1 _06311_ (.A1(\u_glbl_reg.reg_15[2] ),
    .A2(net655),
    .B1(_01823_),
    .X(_01824_));
 sky130_fd_sc_hd__a22o_1 _06312_ (.A1(\u_glbl_reg.reg_16[2] ),
    .A2(net1125),
    .B1(net620),
    .B2(\u_glbl_reg.reg_3[2] ),
    .X(_01825_));
 sky130_fd_sc_hd__a221o_1 _06313_ (.A1(\u_glbl_reg.reg_19[2] ),
    .A2(net641),
    .B1(net607),
    .B2(\u_glbl_reg.cfg_ref_pll_div[2] ),
    .C1(_01825_),
    .X(_01826_));
 sky130_fd_sc_hd__or4_2 _06314_ (.A(_01820_),
    .B(_01822_),
    .C(_01824_),
    .D(_01826_),
    .X(_01827_));
 sky130_fd_sc_hd__nand2_1 _06315_ (.A(\u_glbl_reg.u_random.n1_plus_n0[17] ),
    .B(\u_glbl_reg.u_random.n0[2] ),
    .Y(_01828_));
 sky130_fd_sc_hd__or2_1 _06316_ (.A(\u_glbl_reg.u_random.n1_plus_n0[17] ),
    .B(\u_glbl_reg.u_random.n0[2] ),
    .X(_01829_));
 sky130_fd_sc_hd__nand2_2 _06317_ (.A(_01828_),
    .B(_01829_),
    .Y(_01830_));
 sky130_fd_sc_hd__o21ai_4 _06318_ (.A1(_01790_),
    .A2(_01803_),
    .B1(_01802_),
    .Y(_01831_));
 sky130_fd_sc_hd__xnor2_4 _06319_ (.A(_01830_),
    .B(_01831_),
    .Y(_01832_));
 sky130_fd_sc_hd__a22o_1 _06320_ (.A1(net487),
    .A2(net682),
    .B1(net612),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ),
    .X(_01833_));
 sky130_fd_sc_hd__a221o_1 _06321_ (.A1(\u_glbl_reg.reg_23[2] ),
    .A2(net627),
    .B1(net606),
    .B2(net1098),
    .C1(_01833_),
    .X(_01834_));
 sky130_fd_sc_hd__a221o_1 _06322_ (.A1(net2223),
    .A2(net561),
    .B1(net595),
    .B2(_01832_),
    .C1(_01834_),
    .X(_01835_));
 sky130_fd_sc_hd__or2_1 _06323_ (.A(_01827_),
    .B(_01835_),
    .X(\u_glbl_reg.reg_out[2] ));
 sky130_fd_sc_hd__a21bo_1 _06324_ (.A1(_01829_),
    .A2(_01831_),
    .B1_N(_01828_),
    .X(_01836_));
 sky130_fd_sc_hd__nand2_1 _06325_ (.A(\u_glbl_reg.u_random.n1_plus_n0[18] ),
    .B(\u_glbl_reg.u_random.n0[3] ),
    .Y(_01837_));
 sky130_fd_sc_hd__or2_1 _06326_ (.A(\u_glbl_reg.u_random.n1_plus_n0[18] ),
    .B(\u_glbl_reg.u_random.n0[3] ),
    .X(_01838_));
 sky130_fd_sc_hd__nand3_2 _06327_ (.A(_01836_),
    .B(_01837_),
    .C(_01838_),
    .Y(_01839_));
 sky130_fd_sc_hd__a21o_1 _06328_ (.A1(_01837_),
    .A2(_01838_),
    .B1(_01836_),
    .X(_01840_));
 sky130_fd_sc_hd__a22o_1 _06329_ (.A1(\u_glbl_reg.reg_17[3] ),
    .A2(net649),
    .B1(net646),
    .B2(\u_glbl_reg.reg_18[3] ),
    .X(_01841_));
 sky130_fd_sc_hd__a22o_1 _06330_ (.A1(\u_glbl_reg.reg_19[3] ),
    .A2(net642),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[3] ),
    .X(_01842_));
 sky130_fd_sc_hd__a221o_1 _06331_ (.A1(\u_glbl_reg.reg_3[3] ),
    .A2(net621),
    .B1(net613),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ),
    .C1(_01841_),
    .X(_01843_));
 sky130_fd_sc_hd__a22o_1 _06332_ (.A1(\u_glbl_reg.reg_23[3] ),
    .A2(net625),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[3] ),
    .X(_01844_));
 sky130_fd_sc_hd__a221o_1 _06333_ (.A1(\u_glbl_reg.reg_15[3] ),
    .A2(net655),
    .B1(net589),
    .B2(net184),
    .C1(_01844_),
    .X(_01845_));
 sky130_fd_sc_hd__a22o_1 _06334_ (.A1(net459),
    .A2(net690),
    .B1(net608),
    .B2(net226),
    .X(_01846_));
 sky130_fd_sc_hd__a211o_1 _06335_ (.A1(\u_glbl_reg.cfg_multi_func_sel[3] ),
    .A2(net617),
    .B1(_01843_),
    .C1(_01845_),
    .X(_01847_));
 sky130_fd_sc_hd__a221o_2 _06336_ (.A1(\u_glbl_reg.reg_20[3] ),
    .A2(net638),
    .B1(net634),
    .B2(\u_glbl_reg.reg_21[3] ),
    .C1(_01847_),
    .X(_01848_));
 sky130_fd_sc_hd__a221o_1 _06337_ (.A1(net490),
    .A2(net683),
    .B1(net1124),
    .B2(\u_glbl_reg.reg_16[3] ),
    .C1(_01846_),
    .X(_01849_));
 sky130_fd_sc_hd__a221o_1 _06338_ (.A1(\u_glbl_reg.cfg_rst_ctrl[3] ),
    .A2(net699),
    .B1(net603),
    .B2(net1097),
    .C1(_01842_),
    .X(_01850_));
 sky130_fd_sc_hd__a211o_2 _06339_ (.A1(net2011),
    .A2(net561),
    .B1(_01849_),
    .C1(_01850_),
    .X(_01851_));
 sky130_fd_sc_hd__a31o_1 _06340_ (.A1(net593),
    .A2(_01839_),
    .A3(_01840_),
    .B1(_01851_),
    .X(_01852_));
 sky130_fd_sc_hd__or2_1 _06341_ (.A(_01848_),
    .B(net2012),
    .X(\u_glbl_reg.reg_out[3] ));
 sky130_fd_sc_hd__a21boi_1 _06342_ (.A1(_01836_),
    .A2(_01838_),
    .B1_N(_01837_),
    .Y(_01853_));
 sky130_fd_sc_hd__or2_1 _06343_ (.A(\u_glbl_reg.u_random.n1_plus_n0[19] ),
    .B(\u_glbl_reg.u_random.n0[4] ),
    .X(_01854_));
 sky130_fd_sc_hd__nand2_1 _06344_ (.A(\u_glbl_reg.u_random.n1_plus_n0[19] ),
    .B(\u_glbl_reg.u_random.n0[4] ),
    .Y(_01855_));
 sky130_fd_sc_hd__nand2_1 _06345_ (.A(_01854_),
    .B(_01855_),
    .Y(_01856_));
 sky130_fd_sc_hd__or2_2 _06346_ (.A(_01853_),
    .B(_01856_),
    .X(_01857_));
 sky130_fd_sc_hd__a21oi_2 _06347_ (.A1(_01853_),
    .A2(_01856_),
    .B1(_01789_),
    .Y(_01858_));
 sky130_fd_sc_hd__a22o_1 _06348_ (.A1(\u_glbl_reg.reg_15[4] ),
    .A2(net655),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[4] ),
    .X(_01859_));
 sky130_fd_sc_hd__a221o_2 _06349_ (.A1(\u_glbl_reg.reg_18[4] ),
    .A2(net645),
    .B1(net589),
    .B2(net185),
    .C1(_01859_),
    .X(_01860_));
 sky130_fd_sc_hd__a22o_1 _06350_ (.A1(\u_glbl_reg.reg_19[4] ),
    .A2(net641),
    .B1(net603),
    .B2(net1096),
    .X(_01861_));
 sky130_fd_sc_hd__a221o_1 _06351_ (.A1(\u_glbl_reg.cfg_rst_ctrl[4] ),
    .A2(net698),
    .B1(net612),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ),
    .C1(_01861_),
    .X(_01862_));
 sky130_fd_sc_hd__a22o_1 _06352_ (.A1(\u_glbl_reg.reg_23[4] ),
    .A2(net625),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[4] ),
    .X(_01863_));
 sky130_fd_sc_hd__a221o_1 _06353_ (.A1(net491),
    .A2(net682),
    .B1(net650),
    .B2(\u_glbl_reg.reg_17[4] ),
    .C1(_01863_),
    .X(_01864_));
 sky130_fd_sc_hd__a22o_1 _06354_ (.A1(\u_glbl_reg.reg_16[4] ),
    .A2(net1125),
    .B1(net609),
    .B2(\u_glbl_reg.reg_7[4] ),
    .X(_01865_));
 sky130_fd_sc_hd__a221o_1 _06355_ (.A1(\u_glbl_reg.cfg_mon_sel[0] ),
    .A2(net690),
    .B1(net621),
    .B2(\u_glbl_reg.reg_3[4] ),
    .C1(_01865_),
    .X(_01866_));
 sky130_fd_sc_hd__a211o_1 _06356_ (.A1(\u_glbl_reg.cfg_multi_func_sel[4] ),
    .A2(net617),
    .B1(_01862_),
    .C1(_01864_),
    .X(_01867_));
 sky130_fd_sc_hd__a221o_1 _06357_ (.A1(\u_glbl_reg.reg_20[4] ),
    .A2(net638),
    .B1(net633),
    .B2(\u_glbl_reg.reg_21[4] ),
    .C1(_01867_),
    .X(_01868_));
 sky130_fd_sc_hd__a211o_1 _06358_ (.A1(net1988),
    .A2(net561),
    .B1(_01866_),
    .C1(_01868_),
    .X(_01869_));
 sky130_fd_sc_hd__a211o_1 _06359_ (.A1(_01857_),
    .A2(_01858_),
    .B1(_01860_),
    .C1(_01869_),
    .X(\u_glbl_reg.reg_out[4] ));
 sky130_fd_sc_hd__nand2_1 _06360_ (.A(\u_glbl_reg.u_random.n1_plus_n0[20] ),
    .B(\u_glbl_reg.u_random.n0[5] ),
    .Y(_01870_));
 sky130_fd_sc_hd__or2_1 _06361_ (.A(\u_glbl_reg.u_random.n1_plus_n0[20] ),
    .B(\u_glbl_reg.u_random.n0[5] ),
    .X(_01871_));
 sky130_fd_sc_hd__nand2_1 _06362_ (.A(_01870_),
    .B(_01871_),
    .Y(_01872_));
 sky130_fd_sc_hd__nand2_1 _06363_ (.A(_01855_),
    .B(_01857_),
    .Y(_01873_));
 sky130_fd_sc_hd__a31o_1 _06364_ (.A1(_01870_),
    .A2(_01871_),
    .A3(_01873_),
    .B1(_01789_),
    .X(_01874_));
 sky130_fd_sc_hd__a31oi_4 _06365_ (.A1(_01855_),
    .A2(_01857_),
    .A3(_01872_),
    .B1(_01874_),
    .Y(_01875_));
 sky130_fd_sc_hd__a22o_1 _06366_ (.A1(\u_glbl_reg.cfg_mon_sel[1] ),
    .A2(net686),
    .B1(net625),
    .B2(\u_glbl_reg.reg_23[5] ),
    .X(_01876_));
 sky130_fd_sc_hd__a22o_1 _06367_ (.A1(net492),
    .A2(net682),
    .B1(net642),
    .B2(\u_glbl_reg.reg_19[5] ),
    .X(_01877_));
 sky130_fd_sc_hd__a22o_1 _06368_ (.A1(\u_glbl_reg.reg_18[5] ),
    .A2(net646),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[5] ),
    .X(_01878_));
 sky130_fd_sc_hd__a22o_1 _06369_ (.A1(\u_glbl_reg.cfg_rst_ctrl[5] ),
    .A2(net699),
    .B1(net607),
    .B2(\u_glbl_reg.reg_7[5] ),
    .X(_01879_));
 sky130_fd_sc_hd__a22o_1 _06370_ (.A1(\u_glbl_reg.reg_16[5] ),
    .A2(net1125),
    .B1(net650),
    .B2(\u_glbl_reg.reg_17[5] ),
    .X(_01880_));
 sky130_fd_sc_hd__a211o_1 _06371_ (.A1(net2013),
    .A2(net560),
    .B1(_01879_),
    .C1(_01880_),
    .X(_01881_));
 sky130_fd_sc_hd__a221o_1 _06372_ (.A1(\u_glbl_reg.reg_22[5] ),
    .A2(net629),
    .B1(net604),
    .B2(net1095),
    .C1(_01877_),
    .X(_01882_));
 sky130_fd_sc_hd__a221o_1 _06373_ (.A1(\u_glbl_reg.reg_15[5] ),
    .A2(net655),
    .B1(net589),
    .B2(net186),
    .C1(_01876_),
    .X(_01883_));
 sky130_fd_sc_hd__a221o_1 _06374_ (.A1(\u_glbl_reg.reg_3[5] ),
    .A2(net621),
    .B1(net613),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[5] ),
    .C1(_01878_),
    .X(_01884_));
 sky130_fd_sc_hd__a211o_1 _06375_ (.A1(\u_glbl_reg.cfg_multi_func_sel[5] ),
    .A2(net619),
    .B1(_01883_),
    .C1(_01884_),
    .X(_01885_));
 sky130_fd_sc_hd__a221o_1 _06376_ (.A1(\u_glbl_reg.reg_20[5] ),
    .A2(net638),
    .B1(net634),
    .B2(\u_glbl_reg.reg_21[5] ),
    .C1(_01885_),
    .X(_01886_));
 sky130_fd_sc_hd__or4_2 _06377_ (.A(_01875_),
    .B(_01881_),
    .C(_01882_),
    .D(_01886_),
    .X(\u_glbl_reg.reg_out[5] ));
 sky130_fd_sc_hd__or2_1 _06378_ (.A(\u_glbl_reg.u_random.n1_plus_n0[21] ),
    .B(\u_glbl_reg.u_random.n0[6] ),
    .X(_01887_));
 sky130_fd_sc_hd__nand2_1 _06379_ (.A(\u_glbl_reg.u_random.n1_plus_n0[21] ),
    .B(\u_glbl_reg.u_random.n0[6] ),
    .Y(_01888_));
 sky130_fd_sc_hd__nand2_2 _06380_ (.A(_01887_),
    .B(_01888_),
    .Y(_01889_));
 sky130_fd_sc_hd__and3_1 _06381_ (.A(\u_glbl_reg.u_random.n1_plus_n0[19] ),
    .B(\u_glbl_reg.u_random.n0[4] ),
    .C(_01871_),
    .X(_01890_));
 sky130_fd_sc_hd__a21oi_1 _06382_ (.A1(\u_glbl_reg.u_random.n1_plus_n0[20] ),
    .A2(\u_glbl_reg.u_random.n0[5] ),
    .B1(_01890_),
    .Y(_01891_));
 sky130_fd_sc_hd__o31a_2 _06383_ (.A1(_01853_),
    .A2(_01856_),
    .A3(_01872_),
    .B1(_01891_),
    .X(_01892_));
 sky130_fd_sc_hd__xor2_4 _06384_ (.A(_01889_),
    .B(_01892_),
    .X(_01893_));
 sky130_fd_sc_hd__a22o_1 _06385_ (.A1(\u_glbl_reg.cfg_rtc_clk_ctrl[6] ),
    .A2(net613),
    .B1(net603),
    .B2(net1094),
    .X(_01894_));
 sky130_fd_sc_hd__a22o_1 _06386_ (.A1(\u_glbl_reg.reg_20[6] ),
    .A2(net638),
    .B1(net619),
    .B2(\u_glbl_reg.cfg_multi_func_sel[6] ),
    .X(_01895_));
 sky130_fd_sc_hd__a21o_1 _06387_ (.A1(\u_glbl_reg.reg_21[6] ),
    .A2(net634),
    .B1(_01895_),
    .X(_01896_));
 sky130_fd_sc_hd__a22o_1 _06388_ (.A1(\u_glbl_reg.reg_18[6] ),
    .A2(net645),
    .B1(net608),
    .B2(\u_glbl_reg.reg_7[6] ),
    .X(_01897_));
 sky130_fd_sc_hd__a22o_1 _06389_ (.A1(\u_glbl_reg.reg_22[6] ),
    .A2(net632),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[6] ),
    .X(_01898_));
 sky130_fd_sc_hd__a22o_1 _06390_ (.A1(\u_glbl_reg.reg_16[6] ),
    .A2(net1125),
    .B1(net650),
    .B2(\u_glbl_reg.reg_17[6] ),
    .X(_01899_));
 sky130_fd_sc_hd__a221o_1 _06391_ (.A1(\u_glbl_reg.reg_15[6] ),
    .A2(net656),
    .B1(net642),
    .B2(\u_glbl_reg.reg_19[6] ),
    .C1(_01898_),
    .X(_01900_));
 sky130_fd_sc_hd__a221o_1 _06392_ (.A1(\u_glbl_reg.cfg_rst_ctrl[6] ),
    .A2(net698),
    .B1(net590),
    .B2(net187),
    .C1(_01897_),
    .X(_01901_));
 sky130_fd_sc_hd__a211o_1 _06393_ (.A1(net2091),
    .A2(net561),
    .B1(_01900_),
    .C1(_01901_),
    .X(_01902_));
 sky130_fd_sc_hd__a221o_1 _06394_ (.A1(net493),
    .A2(net683),
    .B1(net621),
    .B2(\u_glbl_reg.reg_3[6] ),
    .C1(_01899_),
    .X(_01903_));
 sky130_fd_sc_hd__a221o_1 _06395_ (.A1(\u_glbl_reg.cfg_mon_sel[2] ),
    .A2(net686),
    .B1(net625),
    .B2(\u_glbl_reg.reg_23[6] ),
    .C1(_01894_),
    .X(_01904_));
 sky130_fd_sc_hd__or3_1 _06396_ (.A(_01896_),
    .B(_01903_),
    .C(_01904_),
    .X(_01905_));
 sky130_fd_sc_hd__a211o_1 _06397_ (.A1(net595),
    .A2(_01893_),
    .B1(_01902_),
    .C1(_01905_),
    .X(\u_glbl_reg.reg_out[6] ));
 sky130_fd_sc_hd__nand2_1 _06398_ (.A(\u_glbl_reg.u_random.n1_plus_n0[22] ),
    .B(\u_glbl_reg.u_random.n0[7] ),
    .Y(_01906_));
 sky130_fd_sc_hd__or2_1 _06399_ (.A(\u_glbl_reg.u_random.n1_plus_n0[22] ),
    .B(\u_glbl_reg.u_random.n0[7] ),
    .X(_01907_));
 sky130_fd_sc_hd__nand2_1 _06400_ (.A(_01906_),
    .B(_01907_),
    .Y(_01908_));
 sky130_fd_sc_hd__o21a_1 _06401_ (.A1(_01889_),
    .A2(_01892_),
    .B1(_01888_),
    .X(_01909_));
 sky130_fd_sc_hd__o21ai_1 _06402_ (.A1(_01908_),
    .A2(_01909_),
    .B1(net594),
    .Y(_01910_));
 sky130_fd_sc_hd__a21oi_4 _06403_ (.A1(_01908_),
    .A2(_01909_),
    .B1(_01910_),
    .Y(_01911_));
 sky130_fd_sc_hd__a22o_1 _06404_ (.A1(net494),
    .A2(net682),
    .B1(net608),
    .B2(\u_glbl_reg.reg_7[7] ),
    .X(_01912_));
 sky130_fd_sc_hd__a22o_1 _06405_ (.A1(\u_glbl_reg.reg_23[7] ),
    .A2(net625),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[7] ),
    .X(_01913_));
 sky130_fd_sc_hd__a22o_1 _06406_ (.A1(\u_glbl_reg.reg_19[7] ),
    .A2(net641),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[7] ),
    .X(_01914_));
 sky130_fd_sc_hd__a22o_1 _06407_ (.A1(\u_glbl_reg.reg_18[7] ),
    .A2(net646),
    .B1(net621),
    .B2(\u_glbl_reg.reg_3[7] ),
    .X(_01915_));
 sky130_fd_sc_hd__a221o_1 _06408_ (.A1(\u_glbl_reg.reg_15[7] ),
    .A2(net655),
    .B1(net589),
    .B2(net188),
    .C1(_01913_),
    .X(_01916_));
 sky130_fd_sc_hd__a221o_1 _06409_ (.A1(\u_glbl_reg.cfg_mon_sel[3] ),
    .A2(net686),
    .B1(net612),
    .B2(\u_glbl_reg.cfg_rtc_clk_ctrl[7] ),
    .C1(_01915_),
    .X(_01917_));
 sky130_fd_sc_hd__a211o_1 _06410_ (.A1(\u_glbl_reg.cfg_multi_func_sel[7] ),
    .A2(net616),
    .B1(_01916_),
    .C1(_01917_),
    .X(_01918_));
 sky130_fd_sc_hd__a221o_1 _06411_ (.A1(\u_glbl_reg.reg_20[7] ),
    .A2(net638),
    .B1(net634),
    .B2(\u_glbl_reg.reg_21[7] ),
    .C1(_01918_),
    .X(_01919_));
 sky130_fd_sc_hd__a221o_1 _06412_ (.A1(\u_glbl_reg.reg_16[7] ),
    .A2(net1124),
    .B1(net650),
    .B2(\u_glbl_reg.reg_17[7] ),
    .C1(_01912_),
    .X(_01920_));
 sky130_fd_sc_hd__a221o_1 _06413_ (.A1(\u_glbl_reg.cfg_rst_ctrl[7] ),
    .A2(net699),
    .B1(net604),
    .B2(net1093),
    .C1(_01914_),
    .X(_01921_));
 sky130_fd_sc_hd__a211o_1 _06414_ (.A1(net2097),
    .A2(net560),
    .B1(_01920_),
    .C1(_01921_),
    .X(_01922_));
 sky130_fd_sc_hd__or3_1 _06415_ (.A(_01911_),
    .B(_01919_),
    .C(net2098),
    .X(\u_glbl_reg.reg_out[7] ));
 sky130_fd_sc_hd__or2_1 _06416_ (.A(\u_glbl_reg.u_random.n1_plus_n0[23] ),
    .B(net1889),
    .X(_01923_));
 sky130_fd_sc_hd__nand2_1 _06417_ (.A(\u_glbl_reg.u_random.n1_plus_n0[23] ),
    .B(net1889),
    .Y(_01924_));
 sky130_fd_sc_hd__nand2_2 _06418_ (.A(_01923_),
    .B(_01924_),
    .Y(_01925_));
 sky130_fd_sc_hd__and3_1 _06419_ (.A(\u_glbl_reg.u_random.n1_plus_n0[21] ),
    .B(\u_glbl_reg.u_random.n0[6] ),
    .C(_01907_),
    .X(_01926_));
 sky130_fd_sc_hd__a21oi_1 _06420_ (.A1(\u_glbl_reg.u_random.n1_plus_n0[22] ),
    .A2(\u_glbl_reg.u_random.n0[7] ),
    .B1(_01926_),
    .Y(_01927_));
 sky130_fd_sc_hd__o31a_2 _06421_ (.A1(_01889_),
    .A2(_01892_),
    .A3(_01908_),
    .B1(_01927_),
    .X(_01928_));
 sky130_fd_sc_hd__nand2_1 _06422_ (.A(_01925_),
    .B(_01928_),
    .Y(_01929_));
 sky130_fd_sc_hd__o21a_1 _06423_ (.A1(_01925_),
    .A2(_01928_),
    .B1(net593),
    .X(_01930_));
 sky130_fd_sc_hd__a22o_1 _06424_ (.A1(\u_glbl_reg.reg_19[8] ),
    .A2(net643),
    .B1(net606),
    .B2(net223),
    .X(_01931_));
 sky130_fd_sc_hd__a22o_1 _06425_ (.A1(\u_glbl_reg.reg_16[8] ),
    .A2(net1128),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[8] ),
    .X(_01932_));
 sky130_fd_sc_hd__a22o_1 _06426_ (.A1(\u_glbl_reg.reg_23[8] ),
    .A2(net627),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[8] ),
    .X(_01933_));
 sky130_fd_sc_hd__a221o_1 _06427_ (.A1(net495),
    .A2(net684),
    .B1(net651),
    .B2(\u_glbl_reg.reg_17[8] ),
    .C1(_01933_),
    .X(_01934_));
 sky130_fd_sc_hd__a221o_1 _06428_ (.A1(\u_glbl_reg.cfg_rst_ctrl[8] ),
    .A2(net700),
    .B1(net614),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[0] ),
    .C1(_01931_),
    .X(_01935_));
 sky130_fd_sc_hd__a22o_1 _06429_ (.A1(\u_glbl_reg.reg_15[8] ),
    .A2(net657),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[8] ),
    .X(_01936_));
 sky130_fd_sc_hd__a221o_1 _06430_ (.A1(\u_glbl_reg.reg_18[8] ),
    .A2(net647),
    .B1(net592),
    .B2(net189),
    .C1(_01936_),
    .X(_01937_));
 sky130_fd_sc_hd__a221o_1 _06431_ (.A1(\u_glbl_reg.cfg_gpio_dgmode ),
    .A2(net688),
    .B1(net623),
    .B2(\u_glbl_reg.reg_3[8] ),
    .C1(_01932_),
    .X(_01938_));
 sky130_fd_sc_hd__a211o_1 _06432_ (.A1(\u_glbl_reg.cfg_multi_func_sel[8] ),
    .A2(net617),
    .B1(_01934_),
    .C1(_01935_),
    .X(_01939_));
 sky130_fd_sc_hd__a221o_1 _06433_ (.A1(\u_glbl_reg.reg_20[8] ),
    .A2(net639),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[8] ),
    .C1(_01939_),
    .X(_01940_));
 sky130_fd_sc_hd__a211o_1 _06434_ (.A1(net1959),
    .A2(net562),
    .B1(_01938_),
    .C1(_01940_),
    .X(_01941_));
 sky130_fd_sc_hd__a211o_1 _06435_ (.A1(_01929_),
    .A2(_01930_),
    .B1(_01937_),
    .C1(net1960),
    .X(\u_glbl_reg.reg_out[8] ));
 sky130_fd_sc_hd__nand2_1 _06436_ (.A(\u_glbl_reg.u_random.n1_plus_n0[24] ),
    .B(net1881),
    .Y(_01942_));
 sky130_fd_sc_hd__or2_1 _06437_ (.A(\u_glbl_reg.u_random.n1_plus_n0[24] ),
    .B(\u_glbl_reg.u_random.n0[9] ),
    .X(_01943_));
 sky130_fd_sc_hd__nand2_1 _06438_ (.A(_01942_),
    .B(_01943_),
    .Y(_01944_));
 sky130_fd_sc_hd__o21ai_1 _06439_ (.A1(_01925_),
    .A2(_01928_),
    .B1(_01924_),
    .Y(_01945_));
 sky130_fd_sc_hd__xnor2_2 _06440_ (.A(_01944_),
    .B(_01945_),
    .Y(_01946_));
 sky130_fd_sc_hd__a22o_1 _06441_ (.A1(\u_glbl_reg.reg_15[9] ),
    .A2(net656),
    .B1(net614),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[1] ),
    .X(_01947_));
 sky130_fd_sc_hd__a221o_1 _06442_ (.A1(\u_glbl_reg.reg_7[9] ),
    .A2(net610),
    .B1(net561),
    .B2(net2031),
    .C1(_01947_),
    .X(_01948_));
 sky130_fd_sc_hd__a221o_1 _06443_ (.A1(\u_glbl_reg.reg_16[9] ),
    .A2(net1131),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[9] ),
    .C1(_01786_),
    .X(_01949_));
 sky130_fd_sc_hd__a221o_1 _06444_ (.A1(\u_glbl_reg.reg_20[9] ),
    .A2(_01550_),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[9] ),
    .C1(_01949_),
    .X(_01950_));
 sky130_fd_sc_hd__a22o_1 _06445_ (.A1(net496),
    .A2(net683),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[9] ),
    .X(_01951_));
 sky130_fd_sc_hd__a221o_1 _06446_ (.A1(\u_glbl_reg.reg_18[9] ),
    .A2(net648),
    .B1(net622),
    .B2(\u_glbl_reg.reg_3[9] ),
    .C1(_01951_),
    .X(_01952_));
 sky130_fd_sc_hd__a22o_1 _06447_ (.A1(\u_glbl_reg.reg_17[9] ),
    .A2(net651),
    .B1(net591),
    .B2(net190),
    .X(_01953_));
 sky130_fd_sc_hd__a221o_1 _06448_ (.A1(\u_glbl_reg.cfg_rst_ctrl[9] ),
    .A2(net700),
    .B1(net642),
    .B2(\u_glbl_reg.reg_19[9] ),
    .C1(_01953_),
    .X(_01954_));
 sky130_fd_sc_hd__a22o_1 _06449_ (.A1(\u_glbl_reg.reg_23[9] ),
    .A2(net627),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[9] ),
    .X(_01955_));
 sky130_fd_sc_hd__a221o_1 _06450_ (.A1(\u_glbl_reg.reg_2[9] ),
    .A2(net687),
    .B1(net604),
    .B2(net224),
    .C1(_01955_),
    .X(_01956_));
 sky130_fd_sc_hd__or2_1 _06451_ (.A(_01954_),
    .B(_01956_),
    .X(_01957_));
 sky130_fd_sc_hd__or4_2 _06452_ (.A(_01948_),
    .B(_01950_),
    .C(_01952_),
    .D(_01957_),
    .X(_01958_));
 sky130_fd_sc_hd__a21o_1 _06453_ (.A1(net593),
    .A2(_01946_),
    .B1(net2032),
    .X(\u_glbl_reg.reg_out[9] ));
 sky130_fd_sc_hd__or2_1 _06454_ (.A(\u_glbl_reg.u_random.n1_plus_n0[25] ),
    .B(\u_glbl_reg.u_random.n0[10] ),
    .X(_01959_));
 sky130_fd_sc_hd__nand2_1 _06455_ (.A(\u_glbl_reg.u_random.n1_plus_n0[25] ),
    .B(\u_glbl_reg.u_random.n0[10] ),
    .Y(_01960_));
 sky130_fd_sc_hd__nand2_1 _06456_ (.A(_01959_),
    .B(_01960_),
    .Y(_01961_));
 sky130_fd_sc_hd__a21bo_1 _06457_ (.A1(_01924_),
    .A2(_01942_),
    .B1_N(_01943_),
    .X(_01962_));
 sky130_fd_sc_hd__or2_1 _06458_ (.A(_01925_),
    .B(_01944_),
    .X(_01963_));
 sky130_fd_sc_hd__or2_1 _06459_ (.A(_01928_),
    .B(_01963_),
    .X(_01964_));
 sky130_fd_sc_hd__a21o_1 _06460_ (.A1(_01962_),
    .A2(_01964_),
    .B1(_01961_),
    .X(_01965_));
 sky130_fd_sc_hd__nand2_1 _06461_ (.A(net594),
    .B(_01965_),
    .Y(_01966_));
 sky130_fd_sc_hd__a31o_1 _06462_ (.A1(_01961_),
    .A2(_01962_),
    .A3(_01964_),
    .B1(_01966_),
    .X(_01967_));
 sky130_fd_sc_hd__a22o_1 _06463_ (.A1(\u_glbl_reg.reg_21[10] ),
    .A2(net636),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .X(_01968_));
 sky130_fd_sc_hd__a221o_1 _06464_ (.A1(\u_glbl_reg.reg_20[10] ),
    .A2(net639),
    .B1(net627),
    .B2(\u_glbl_reg.reg_23[10] ),
    .C1(_01786_),
    .X(_01969_));
 sky130_fd_sc_hd__or2_1 _06465_ (.A(_01968_),
    .B(_01969_),
    .X(_01970_));
 sky130_fd_sc_hd__a22o_1 _06466_ (.A1(\u_glbl_reg.reg_16[10] ),
    .A2(net1128),
    .B1(net652),
    .B2(\u_glbl_reg.reg_17[10] ),
    .X(_01971_));
 sky130_fd_sc_hd__a221o_1 _06467_ (.A1(\u_glbl_reg.cfg_rst_ctrl[10] ),
    .A2(net700),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[10] ),
    .C1(_01971_),
    .X(_01972_));
 sky130_fd_sc_hd__a22o_1 _06468_ (.A1(net200),
    .A2(net604),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[10] ),
    .X(_01973_));
 sky130_fd_sc_hd__a221o_1 _06469_ (.A1(\u_glbl_reg.reg_7[10] ),
    .A2(net610),
    .B1(net561),
    .B2(net2050),
    .C1(_01973_),
    .X(_01974_));
 sky130_fd_sc_hd__a22o_1 _06470_ (.A1(\u_glbl_reg.reg_19[10] ),
    .A2(net642),
    .B1(net591),
    .B2(net160),
    .X(_01975_));
 sky130_fd_sc_hd__a221o_1 _06471_ (.A1(net466),
    .A2(net684),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[10] ),
    .C1(_01975_),
    .X(_01976_));
 sky130_fd_sc_hd__a22o_1 _06472_ (.A1(\u_glbl_reg.reg_15[10] ),
    .A2(net656),
    .B1(net622),
    .B2(\u_glbl_reg.reg_3[10] ),
    .X(_01977_));
 sky130_fd_sc_hd__a22o_1 _06473_ (.A1(\u_glbl_reg.reg_2[10] ),
    .A2(net687),
    .B1(net614),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[2] ),
    .X(_01978_));
 sky130_fd_sc_hd__or4_2 _06474_ (.A(_01974_),
    .B(_01976_),
    .C(_01977_),
    .D(_01978_),
    .X(_01979_));
 sky130_fd_sc_hd__or4b_1 _06475_ (.A(_01970_),
    .B(_01972_),
    .C(net2051),
    .D_N(_01967_),
    .X(\u_glbl_reg.reg_out[10] ));
 sky130_fd_sc_hd__and2_1 _06476_ (.A(\u_glbl_reg.u_random.n1_plus_n0[26] ),
    .B(\u_glbl_reg.u_random.n0[11] ),
    .X(_01980_));
 sky130_fd_sc_hd__nor2_1 _06477_ (.A(\u_glbl_reg.u_random.n1_plus_n0[26] ),
    .B(\u_glbl_reg.u_random.n0[11] ),
    .Y(_01981_));
 sky130_fd_sc_hd__or2_1 _06478_ (.A(_01980_),
    .B(_01981_),
    .X(_01982_));
 sky130_fd_sc_hd__nand2_1 _06479_ (.A(_01960_),
    .B(_01965_),
    .Y(_01983_));
 sky130_fd_sc_hd__xnor2_2 _06480_ (.A(_01982_),
    .B(_01983_),
    .Y(_01984_));
 sky130_fd_sc_hd__a22o_1 _06481_ (.A1(\u_glbl_reg.reg_19[11] ),
    .A2(net643),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[11] ),
    .X(_01985_));
 sky130_fd_sc_hd__a22o_1 _06482_ (.A1(\u_glbl_reg.reg_17[11] ),
    .A2(net651),
    .B1(net648),
    .B2(\u_glbl_reg.reg_18[11] ),
    .X(_01986_));
 sky130_fd_sc_hd__a221o_1 _06483_ (.A1(\u_glbl_reg.reg_3[11] ),
    .A2(net622),
    .B1(net614),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[3] ),
    .C1(_01986_),
    .X(_01987_));
 sky130_fd_sc_hd__a221o_1 _06484_ (.A1(\u_glbl_reg.cfg_rst_ctrl[11] ),
    .A2(net700),
    .B1(net604),
    .B2(net201),
    .C1(_01985_),
    .X(_01988_));
 sky130_fd_sc_hd__a22o_1 _06485_ (.A1(\u_glbl_reg.reg_2[11] ),
    .A2(net687),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[11] ),
    .X(_01989_));
 sky130_fd_sc_hd__a221o_1 _06486_ (.A1(net467),
    .A2(_01146_),
    .B1(net1128),
    .B2(\u_glbl_reg.reg_16[11] ),
    .C1(_01989_),
    .X(_01990_));
 sky130_fd_sc_hd__a22o_1 _06487_ (.A1(\u_glbl_reg.reg_23[11] ),
    .A2(net627),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[11] ),
    .X(_01991_));
 sky130_fd_sc_hd__a221o_1 _06488_ (.A1(\u_glbl_reg.reg_15[11] ),
    .A2(net656),
    .B1(net591),
    .B2(net161),
    .C1(_01991_),
    .X(_01992_));
 sky130_fd_sc_hd__a211o_1 _06489_ (.A1(net1982),
    .A2(net562),
    .B1(_01988_),
    .C1(_01990_),
    .X(_01993_));
 sky130_fd_sc_hd__a211o_1 _06490_ (.A1(\u_glbl_reg.cfg_multi_func_sel[11] ),
    .A2(net619),
    .B1(_01987_),
    .C1(_01992_),
    .X(_01994_));
 sky130_fd_sc_hd__a221o_1 _06491_ (.A1(\u_glbl_reg.reg_20[11] ),
    .A2(net639),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[11] ),
    .C1(_01994_),
    .X(_01995_));
 sky130_fd_sc_hd__a211o_1 _06492_ (.A1(net595),
    .A2(_01984_),
    .B1(_01993_),
    .C1(_01995_),
    .X(\u_glbl_reg.reg_out[11] ));
 sky130_fd_sc_hd__or2_1 _06493_ (.A(\u_glbl_reg.u_random.n1_plus_n0[27] ),
    .B(\u_glbl_reg.u_random.n0[12] ),
    .X(_01996_));
 sky130_fd_sc_hd__nand2_1 _06494_ (.A(\u_glbl_reg.u_random.n1_plus_n0[27] ),
    .B(\u_glbl_reg.u_random.n0[12] ),
    .Y(_01997_));
 sky130_fd_sc_hd__nand2_1 _06495_ (.A(_01996_),
    .B(_01997_),
    .Y(_01998_));
 sky130_fd_sc_hd__or2_1 _06496_ (.A(_01961_),
    .B(_01982_),
    .X(_01999_));
 sky130_fd_sc_hd__o21ba_1 _06497_ (.A1(_01960_),
    .A2(_01981_),
    .B1_N(_01980_),
    .X(_02000_));
 sky130_fd_sc_hd__o21a_1 _06498_ (.A1(_01962_),
    .A2(_01999_),
    .B1(_02000_),
    .X(_02001_));
 sky130_fd_sc_hd__or2_1 _06499_ (.A(_01963_),
    .B(_01999_),
    .X(_02002_));
 sky130_fd_sc_hd__o21ai_2 _06500_ (.A1(_01928_),
    .A2(_02002_),
    .B1(_02001_),
    .Y(_02003_));
 sky130_fd_sc_hd__xnor2_2 _06501_ (.A(_01998_),
    .B(_02003_),
    .Y(_02004_));
 sky130_fd_sc_hd__a22o_1 _06502_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[4] ),
    .A2(net613),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[12] ),
    .X(_02005_));
 sky130_fd_sc_hd__a211o_1 _06503_ (.A1(\u_glbl_reg.reg_3[12] ),
    .A2(net621),
    .B1(_01786_),
    .C1(_02005_),
    .X(_02006_));
 sky130_fd_sc_hd__a22o_1 _06504_ (.A1(\u_glbl_reg.reg_20[12] ),
    .A2(net638),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[12] ),
    .X(_02007_));
 sky130_fd_sc_hd__a221o_1 _06505_ (.A1(\u_glbl_reg.reg_15[12] ),
    .A2(net657),
    .B1(net644),
    .B2(\u_glbl_reg.reg_19[12] ),
    .C1(_02007_),
    .X(_02008_));
 sky130_fd_sc_hd__a22o_1 _06506_ (.A1(\u_glbl_reg.cfg_rst_ctrl[12] ),
    .A2(net700),
    .B1(net1126),
    .B2(\u_glbl_reg.reg_16[12] ),
    .X(_02009_));
 sky130_fd_sc_hd__a221o_1 _06507_ (.A1(\u_glbl_reg.cfg_multi_func_sel[12] ),
    .A2(net618),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[12] ),
    .C1(_02009_),
    .X(_02010_));
 sky130_fd_sc_hd__a22o_1 _06508_ (.A1(\u_glbl_reg.reg_23[12] ),
    .A2(net627),
    .B1(net591),
    .B2(net162),
    .X(_02011_));
 sky130_fd_sc_hd__a221o_1 _06509_ (.A1(\u_glbl_reg.reg_2[12] ),
    .A2(net687),
    .B1(net684),
    .B2(net468),
    .C1(_02011_),
    .X(_02012_));
 sky130_fd_sc_hd__a22o_1 _06510_ (.A1(\u_glbl_reg.reg_18[12] ),
    .A2(net648),
    .B1(net605),
    .B2(net202),
    .X(_02013_));
 sky130_fd_sc_hd__a221o_1 _06511_ (.A1(\u_glbl_reg.reg_17[12] ),
    .A2(net652),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[12] ),
    .C1(_02013_),
    .X(_02014_));
 sky130_fd_sc_hd__or4_1 _06512_ (.A(_02008_),
    .B(_02010_),
    .C(_02012_),
    .D(_02014_),
    .X(_02015_));
 sky130_fd_sc_hd__a211o_1 _06513_ (.A1(net1990),
    .A2(net561),
    .B1(_02006_),
    .C1(_02015_),
    .X(_02016_));
 sky130_fd_sc_hd__a21o_1 _06514_ (.A1(net595),
    .A2(_02004_),
    .B1(net1991),
    .X(\u_glbl_reg.reg_out[12] ));
 sky130_fd_sc_hd__nand2_1 _06515_ (.A(\u_glbl_reg.u_random.n1_plus_n0[28] ),
    .B(\u_glbl_reg.u_random.n0[13] ),
    .Y(_02017_));
 sky130_fd_sc_hd__nor2_1 _06516_ (.A(\u_glbl_reg.u_random.n1_plus_n0[28] ),
    .B(\u_glbl_reg.u_random.n0[13] ),
    .Y(_02018_));
 sky130_fd_sc_hd__or2_1 _06517_ (.A(\u_glbl_reg.u_random.n1_plus_n0[28] ),
    .B(\u_glbl_reg.u_random.n0[13] ),
    .X(_02019_));
 sky130_fd_sc_hd__nand2_1 _06518_ (.A(_02017_),
    .B(_02019_),
    .Y(_02020_));
 sky130_fd_sc_hd__a21boi_2 _06519_ (.A1(_01996_),
    .A2(_02003_),
    .B1_N(_01997_),
    .Y(_02021_));
 sky130_fd_sc_hd__o21ai_1 _06520_ (.A1(_02020_),
    .A2(_02021_),
    .B1(net594),
    .Y(_02022_));
 sky130_fd_sc_hd__a21oi_4 _06521_ (.A1(_02020_),
    .A2(_02021_),
    .B1(_02022_),
    .Y(_02023_));
 sky130_fd_sc_hd__a22o_1 _06522_ (.A1(\u_glbl_reg.reg_2[13] ),
    .A2(net688),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[13] ),
    .X(_02024_));
 sky130_fd_sc_hd__a22o_1 _06523_ (.A1(net469),
    .A2(net683),
    .B1(net656),
    .B2(\u_glbl_reg.reg_15[13] ),
    .X(_02025_));
 sky130_fd_sc_hd__a22o_1 _06524_ (.A1(\u_glbl_reg.reg_19[13] ),
    .A2(net643),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[13] ),
    .X(_02026_));
 sky130_fd_sc_hd__a22o_1 _06525_ (.A1(\u_glbl_reg.reg_17[13] ),
    .A2(net651),
    .B1(net648),
    .B2(\u_glbl_reg.reg_18[13] ),
    .X(_02027_));
 sky130_fd_sc_hd__a221o_1 _06526_ (.A1(\u_glbl_reg.reg_23[13] ),
    .A2(net627),
    .B1(net591),
    .B2(net163),
    .C1(_02025_),
    .X(_02028_));
 sky130_fd_sc_hd__a221o_1 _06527_ (.A1(\u_glbl_reg.reg_3[13] ),
    .A2(net622),
    .B1(net613),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[5] ),
    .C1(_02027_),
    .X(_02029_));
 sky130_fd_sc_hd__a211o_1 _06528_ (.A1(\u_glbl_reg.cfg_multi_func_sel[13] ),
    .A2(net617),
    .B1(_02028_),
    .C1(_02029_),
    .X(_02030_));
 sky130_fd_sc_hd__a221o_1 _06529_ (.A1(\u_glbl_reg.reg_20[13] ),
    .A2(net639),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[13] ),
    .C1(_02030_),
    .X(_02031_));
 sky130_fd_sc_hd__a221o_1 _06530_ (.A1(\u_glbl_reg.reg_16[13] ),
    .A2(net1128),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[13] ),
    .C1(_02024_),
    .X(_02032_));
 sky130_fd_sc_hd__a221o_1 _06531_ (.A1(\u_glbl_reg.cfg_rst_ctrl[13] ),
    .A2(net700),
    .B1(net606),
    .B2(net203),
    .C1(_02026_),
    .X(_02033_));
 sky130_fd_sc_hd__a211o_1 _06532_ (.A1(net1965),
    .A2(net562),
    .B1(_02032_),
    .C1(_02033_),
    .X(_02034_));
 sky130_fd_sc_hd__or3_1 _06533_ (.A(_02023_),
    .B(_02031_),
    .C(_02034_),
    .X(\u_glbl_reg.reg_out[13] ));
 sky130_fd_sc_hd__or2_1 _06534_ (.A(\u_glbl_reg.u_random.n1_plus_n0[29] ),
    .B(net1909),
    .X(_02035_));
 sky130_fd_sc_hd__nand2_1 _06535_ (.A(\u_glbl_reg.u_random.n1_plus_n0[29] ),
    .B(\u_glbl_reg.u_random.n0[14] ),
    .Y(_02036_));
 sky130_fd_sc_hd__nand2_1 _06536_ (.A(_02035_),
    .B(_02036_),
    .Y(_02037_));
 sky130_fd_sc_hd__a21o_1 _06537_ (.A1(_02017_),
    .A2(_02021_),
    .B1(_02018_),
    .X(_02038_));
 sky130_fd_sc_hd__nand2_1 _06538_ (.A(_02037_),
    .B(_02038_),
    .Y(_02039_));
 sky130_fd_sc_hd__or2_2 _06539_ (.A(_02037_),
    .B(_02038_),
    .X(_02040_));
 sky130_fd_sc_hd__a22o_1 _06540_ (.A1(\u_glbl_reg.reg_22[14] ),
    .A2(net630),
    .B1(net626),
    .B2(\u_glbl_reg.reg_23[14] ),
    .X(_02041_));
 sky130_fd_sc_hd__a22o_1 _06541_ (.A1(\u_glbl_reg.reg_2[14] ),
    .A2(net688),
    .B1(net609),
    .B2(\u_glbl_reg.reg_7[14] ),
    .X(_02042_));
 sky130_fd_sc_hd__a22o_2 _06542_ (.A1(net470),
    .A2(net681),
    .B1(net596),
    .B2(\u_glbl_reg.reg_12[14] ),
    .X(_02043_));
 sky130_fd_sc_hd__a221o_1 _06543_ (.A1(\u_glbl_reg.reg_19[14] ),
    .A2(net643),
    .B1(net623),
    .B2(\u_glbl_reg.reg_3[14] ),
    .C1(_02043_),
    .X(_02044_));
 sky130_fd_sc_hd__a22o_1 _06544_ (.A1(\u_glbl_reg.reg_16[14] ),
    .A2(net1127),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[14] ),
    .X(_02045_));
 sky130_fd_sc_hd__a221o_1 _06545_ (.A1(\u_glbl_reg.cfg_rst_ctrl[14] ),
    .A2(net701),
    .B1(net652),
    .B2(\u_glbl_reg.reg_17[14] ),
    .C1(_02045_),
    .X(_02046_));
 sky130_fd_sc_hd__a221o_1 _06546_ (.A1(\u_glbl_reg.reg_15[14] ),
    .A2(net657),
    .B1(net604),
    .B2(net204),
    .C1(_02041_),
    .X(_02047_));
 sky130_fd_sc_hd__a221o_1 _06547_ (.A1(\u_glbl_reg.cfg_usb_clk_ctrl[6] ),
    .A2(net614),
    .B1(net591),
    .B2(net164),
    .C1(_02042_),
    .X(_02048_));
 sky130_fd_sc_hd__a211o_1 _06548_ (.A1(\u_glbl_reg.cfg_multi_func_sel[14] ),
    .A2(net618),
    .B1(_02047_),
    .C1(_02048_),
    .X(_02049_));
 sky130_fd_sc_hd__a221o_1 _06549_ (.A1(\u_glbl_reg.reg_20[14] ),
    .A2(net639),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[14] ),
    .C1(_02049_),
    .X(_02050_));
 sky130_fd_sc_hd__a211o_1 _06550_ (.A1(net1993),
    .A2(net562),
    .B1(_02044_),
    .C1(_02050_),
    .X(_02051_));
 sky130_fd_sc_hd__a311o_1 _06551_ (.A1(net593),
    .A2(_02039_),
    .A3(_02040_),
    .B1(_02046_),
    .C1(_02051_),
    .X(\u_glbl_reg.reg_out[14] ));
 sky130_fd_sc_hd__or2_1 _06552_ (.A(\u_glbl_reg.u_random.n1_plus_n0[30] ),
    .B(\u_glbl_reg.u_random.n0[15] ),
    .X(_02052_));
 sky130_fd_sc_hd__nand2_1 _06553_ (.A(\u_glbl_reg.u_random.n1_plus_n0[30] ),
    .B(\u_glbl_reg.u_random.n0[15] ),
    .Y(_02053_));
 sky130_fd_sc_hd__nand2_1 _06554_ (.A(_02052_),
    .B(_02053_),
    .Y(_02054_));
 sky130_fd_sc_hd__a21oi_1 _06555_ (.A1(_02036_),
    .A2(_02040_),
    .B1(_02054_),
    .Y(_02055_));
 sky130_fd_sc_hd__a31o_1 _06556_ (.A1(_02036_),
    .A2(_02040_),
    .A3(_02054_),
    .B1(_01789_),
    .X(_02056_));
 sky130_fd_sc_hd__nor2_2 _06557_ (.A(_02055_),
    .B(_02056_),
    .Y(_02057_));
 sky130_fd_sc_hd__a22o_1 _06558_ (.A1(\u_glbl_reg.reg_23[15] ),
    .A2(net627),
    .B1(net597),
    .B2(\u_glbl_reg.reg_12[15] ),
    .X(_02058_));
 sky130_fd_sc_hd__a22o_1 _06559_ (.A1(\u_glbl_reg.reg_2[15] ),
    .A2(net688),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[15] ),
    .X(_02059_));
 sky130_fd_sc_hd__a221o_1 _06560_ (.A1(net471),
    .A2(_01146_),
    .B1(net1128),
    .B2(\u_glbl_reg.reg_16[15] ),
    .C1(_02059_),
    .X(_02060_));
 sky130_fd_sc_hd__a22o_1 _06561_ (.A1(\u_glbl_reg.reg_17[15] ),
    .A2(net651),
    .B1(net648),
    .B2(\u_glbl_reg.reg_18[15] ),
    .X(_02061_));
 sky130_fd_sc_hd__a22o_1 _06562_ (.A1(\u_glbl_reg.reg_19[15] ),
    .A2(net643),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[15] ),
    .X(_02062_));
 sky130_fd_sc_hd__a221o_1 _06563_ (.A1(\u_glbl_reg.cfg_rst_ctrl[15] ),
    .A2(net701),
    .B1(net606),
    .B2(net205),
    .C1(_02062_),
    .X(_02063_));
 sky130_fd_sc_hd__a211o_1 _06564_ (.A1(net1967),
    .A2(net562),
    .B1(_02060_),
    .C1(_02063_),
    .X(_02064_));
 sky130_fd_sc_hd__a221o_1 _06565_ (.A1(\u_glbl_reg.reg_15[15] ),
    .A2(net656),
    .B1(net591),
    .B2(net165),
    .C1(_02058_),
    .X(_02065_));
 sky130_fd_sc_hd__a221o_1 _06566_ (.A1(\u_glbl_reg.reg_3[15] ),
    .A2(net622),
    .B1(net615),
    .B2(\u_glbl_reg.cfg_usb_clk_ctrl[7] ),
    .C1(_02061_),
    .X(_02066_));
 sky130_fd_sc_hd__a211o_1 _06567_ (.A1(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .A2(net617),
    .B1(_02065_),
    .C1(_02066_),
    .X(_02067_));
 sky130_fd_sc_hd__a221o_1 _06568_ (.A1(\u_glbl_reg.reg_20[15] ),
    .A2(net639),
    .B1(net636),
    .B2(\u_glbl_reg.reg_21[15] ),
    .C1(_02067_),
    .X(_02068_));
 sky130_fd_sc_hd__or3_1 _06569_ (.A(_02057_),
    .B(net1968),
    .C(_02068_),
    .X(\u_glbl_reg.reg_out[15] ));
 sky130_fd_sc_hd__or2_1 _06570_ (.A(_02037_),
    .B(_02054_),
    .X(_02069_));
 sky130_fd_sc_hd__or3_1 _06571_ (.A(_01998_),
    .B(_02020_),
    .C(_02069_),
    .X(_02070_));
 sky130_fd_sc_hd__a21bo_1 _06572_ (.A1(_02036_),
    .A2(_02053_),
    .B1_N(_02052_),
    .X(_02071_));
 sky130_fd_sc_hd__o21a_1 _06573_ (.A1(_01997_),
    .A2(_02018_),
    .B1(_02017_),
    .X(_02072_));
 sky130_fd_sc_hd__o221a_1 _06574_ (.A1(_02001_),
    .A2(_02070_),
    .B1(_02072_),
    .B2(_02069_),
    .C1(_02071_),
    .X(_02073_));
 sky130_fd_sc_hd__o31a_2 _06575_ (.A1(_01928_),
    .A2(_02002_),
    .A3(_02070_),
    .B1(_02073_),
    .X(_02074_));
 sky130_fd_sc_hd__or2_1 _06576_ (.A(net2028),
    .B(net1917),
    .X(_02075_));
 sky130_fd_sc_hd__nand2_1 _06577_ (.A(net2028),
    .B(\u_glbl_reg.u_random.n0[16] ),
    .Y(_02076_));
 sky130_fd_sc_hd__nand2_1 _06578_ (.A(_02075_),
    .B(_02076_),
    .Y(_02077_));
 sky130_fd_sc_hd__or2_1 _06579_ (.A(_02074_),
    .B(_02077_),
    .X(_02078_));
 sky130_fd_sc_hd__nand2_1 _06580_ (.A(_02074_),
    .B(_02077_),
    .Y(_02079_));
 sky130_fd_sc_hd__a22o_1 _06581_ (.A1(\u_glbl_reg.reg_20[16] ),
    .A2(net640),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[16] ),
    .X(_02080_));
 sky130_fd_sc_hd__a221o_1 _06582_ (.A1(\u_glbl_reg.reg_2[16] ),
    .A2(net689),
    .B1(net635),
    .B2(\u_glbl_reg.reg_21[16] ),
    .C1(_02080_),
    .X(_02081_));
 sky130_fd_sc_hd__a22o_1 _06583_ (.A1(\u_glbl_reg.reg_23[16] ),
    .A2(net626),
    .B1(net614),
    .B2(\u_glbl_reg.reg_6[16] ),
    .X(_02082_));
 sky130_fd_sc_hd__a211o_1 _06584_ (.A1(net2066),
    .A2(net563),
    .B1(_02081_),
    .C1(_02082_),
    .X(_02083_));
 sky130_fd_sc_hd__a22o_1 _06585_ (.A1(net472),
    .A2(net684),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[16] ),
    .X(_02084_));
 sky130_fd_sc_hd__a221o_1 _06586_ (.A1(\u_glbl_reg.reg_3[16] ),
    .A2(net623),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[16] ),
    .C1(_02084_),
    .X(_02085_));
 sky130_fd_sc_hd__a22o_1 _06587_ (.A1(\u_glbl_reg.reg_15[16] ),
    .A2(net657),
    .B1(net1127),
    .B2(\u_glbl_reg.reg_16[16] ),
    .X(_02086_));
 sky130_fd_sc_hd__a22o_1 _06588_ (.A1(\u_glbl_reg.reg_18[16] ),
    .A2(net647),
    .B1(net605),
    .B2(net206),
    .X(_02087_));
 sky130_fd_sc_hd__a22o_1 _06589_ (.A1(\u_glbl_reg.reg_17[16] ),
    .A2(net652),
    .B1(net592),
    .B2(net166),
    .X(_02088_));
 sky130_fd_sc_hd__a221o_1 _06590_ (.A1(\u_glbl_reg.cfg_rst_ctrl[16] ),
    .A2(net701),
    .B1(net643),
    .B2(\u_glbl_reg.reg_19[16] ),
    .C1(_02088_),
    .X(_02089_));
 sky130_fd_sc_hd__or4_1 _06591_ (.A(_02085_),
    .B(_02086_),
    .C(_02087_),
    .D(_02089_),
    .X(_02090_));
 sky130_fd_sc_hd__or2_1 _06592_ (.A(_02083_),
    .B(_02090_),
    .X(_02091_));
 sky130_fd_sc_hd__a31o_1 _06593_ (.A1(net594),
    .A2(_02078_),
    .A3(_02079_),
    .B1(_02091_),
    .X(\u_glbl_reg.reg_out[16] ));
 sky130_fd_sc_hd__nand2_1 _06594_ (.A(net2008),
    .B(net1884),
    .Y(_02092_));
 sky130_fd_sc_hd__or2_1 _06595_ (.A(net2008),
    .B(\u_glbl_reg.u_random.n0[17] ),
    .X(_02093_));
 sky130_fd_sc_hd__nand2_1 _06596_ (.A(_02092_),
    .B(_02093_),
    .Y(_02094_));
 sky130_fd_sc_hd__o21ai_1 _06597_ (.A1(_02074_),
    .A2(_02077_),
    .B1(net2029),
    .Y(_02095_));
 sky130_fd_sc_hd__xnor2_1 _06598_ (.A(_02094_),
    .B(_02095_),
    .Y(_02096_));
 sky130_fd_sc_hd__a22o_1 _06599_ (.A1(\u_glbl_reg.reg_3[17] ),
    .A2(net623),
    .B1(net605),
    .B2(net207),
    .X(_02097_));
 sky130_fd_sc_hd__a221o_1 _06600_ (.A1(\u_glbl_reg.reg_15[17] ),
    .A2(net657),
    .B1(net562),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ),
    .C1(_02097_),
    .X(_02098_));
 sky130_fd_sc_hd__a22o_1 _06601_ (.A1(\u_glbl_reg.reg_20[17] ),
    .A2(net639),
    .B1(net635),
    .B2(\u_glbl_reg.reg_21[17] ),
    .X(_02099_));
 sky130_fd_sc_hd__a22o_1 _06602_ (.A1(\u_glbl_reg.cfg_rst_ctrl[17] ),
    .A2(net701),
    .B1(net687),
    .B2(\u_glbl_reg.reg_2[17] ),
    .X(_02100_));
 sky130_fd_sc_hd__a221o_1 _06603_ (.A1(\u_glbl_reg.reg_6[17] ),
    .A2(net614),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[17] ),
    .C1(_02100_),
    .X(_02101_));
 sky130_fd_sc_hd__a2111o_1 _06604_ (.A1(\u_glbl_reg.cfg_multi_func_sel[17] ),
    .A2(net619),
    .B1(_02098_),
    .C1(_02099_),
    .D1(_02101_),
    .X(_02102_));
 sky130_fd_sc_hd__a22o_1 _06605_ (.A1(\u_glbl_reg.reg_16[17] ),
    .A2(net1127),
    .B1(net653),
    .B2(\u_glbl_reg.reg_17[17] ),
    .X(_02103_));
 sky130_fd_sc_hd__a22o_1 _06606_ (.A1(\u_glbl_reg.reg_19[17] ),
    .A2(net644),
    .B1(net631),
    .B2(\u_glbl_reg.reg_22[17] ),
    .X(_02104_));
 sky130_fd_sc_hd__a22o_2 _06607_ (.A1(net473),
    .A2(net681),
    .B1(net589),
    .B2(net167),
    .X(_02105_));
 sky130_fd_sc_hd__a221o_1 _06608_ (.A1(\u_glbl_reg.reg_18[17] ),
    .A2(net648),
    .B1(net626),
    .B2(\u_glbl_reg.reg_23[17] ),
    .C1(_02105_),
    .X(_02106_));
 sky130_fd_sc_hd__or4_1 _06609_ (.A(_02102_),
    .B(_02103_),
    .C(_02104_),
    .D(_02106_),
    .X(_02107_));
 sky130_fd_sc_hd__a21o_1 _06610_ (.A1(net593),
    .A2(net2030),
    .B1(_02107_),
    .X(\u_glbl_reg.reg_out[17] ));
 sky130_fd_sc_hd__or2_1 _06611_ (.A(net1984),
    .B(net1931),
    .X(_02108_));
 sky130_fd_sc_hd__nand2_1 _06612_ (.A(net1984),
    .B(net1931),
    .Y(_02109_));
 sky130_fd_sc_hd__nand2_1 _06613_ (.A(_02108_),
    .B(_02109_),
    .Y(_02110_));
 sky130_fd_sc_hd__a21bo_1 _06614_ (.A1(_02076_),
    .A2(_02092_),
    .B1_N(_02093_),
    .X(_02111_));
 sky130_fd_sc_hd__or2_1 _06615_ (.A(_02077_),
    .B(_02094_),
    .X(_02112_));
 sky130_fd_sc_hd__or2_1 _06616_ (.A(_02074_),
    .B(_02112_),
    .X(_02113_));
 sky130_fd_sc_hd__a21o_1 _06617_ (.A1(_02111_),
    .A2(_02113_),
    .B1(_02110_),
    .X(_02114_));
 sky130_fd_sc_hd__nand3_1 _06618_ (.A(_02110_),
    .B(net2009),
    .C(_02113_),
    .Y(_02115_));
 sky130_fd_sc_hd__a22o_1 _06619_ (.A1(\u_glbl_reg.reg_3[18] ),
    .A2(net623),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[18] ),
    .X(_02116_));
 sky130_fd_sc_hd__a221o_1 _06620_ (.A1(\u_glbl_reg.reg_6[18] ),
    .A2(net615),
    .B1(net605),
    .B2(net208),
    .C1(_02116_),
    .X(_02117_));
 sky130_fd_sc_hd__a22o_1 _06621_ (.A1(\u_glbl_reg.reg_23[18] ),
    .A2(net626),
    .B1(net591),
    .B2(net168),
    .X(_02118_));
 sky130_fd_sc_hd__a221o_1 _06622_ (.A1(\u_glbl_reg.cfg_rst_ctrl[18] ),
    .A2(net700),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[18] ),
    .C1(_02118_),
    .X(_02119_));
 sky130_fd_sc_hd__a22o_1 _06623_ (.A1(net474),
    .A2(net684),
    .B1(net1127),
    .B2(\u_glbl_reg.reg_16[18] ),
    .X(_02120_));
 sky130_fd_sc_hd__a221o_1 _06624_ (.A1(\u_glbl_reg.reg_17[18] ),
    .A2(net652),
    .B1(net563),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ),
    .C1(_02120_),
    .X(_02121_));
 sky130_fd_sc_hd__a22o_1 _06625_ (.A1(\u_glbl_reg.reg_19[18] ),
    .A2(net643),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[18] ),
    .X(_02122_));
 sky130_fd_sc_hd__a221o_1 _06626_ (.A1(\u_glbl_reg.reg_2[18] ),
    .A2(net689),
    .B1(net657),
    .B2(\u_glbl_reg.reg_15[18] ),
    .C1(_02122_),
    .X(_02123_));
 sky130_fd_sc_hd__a22o_1 _06627_ (.A1(\u_glbl_reg.reg_21[18] ),
    .A2(net635),
    .B1(net619),
    .B2(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .X(_02124_));
 sky130_fd_sc_hd__a2111o_1 _06628_ (.A1(\u_glbl_reg.reg_20[18] ),
    .A2(net639),
    .B1(_02121_),
    .C1(_02123_),
    .D1(_02124_),
    .X(_02125_));
 sky130_fd_sc_hd__or3_1 _06629_ (.A(_02117_),
    .B(_02119_),
    .C(_02125_),
    .X(_02126_));
 sky130_fd_sc_hd__a31o_1 _06630_ (.A1(net594),
    .A2(_02114_),
    .A3(_02115_),
    .B1(_02126_),
    .X(\u_glbl_reg.reg_out[18] ));
 sky130_fd_sc_hd__and2_1 _06631_ (.A(\u_glbl_reg.u_random.n1_plus_n0[2] ),
    .B(net1927),
    .X(_02127_));
 sky130_fd_sc_hd__nor2_1 _06632_ (.A(\u_glbl_reg.u_random.n1_plus_n0[2] ),
    .B(\u_glbl_reg.u_random.n0[19] ),
    .Y(_02128_));
 sky130_fd_sc_hd__or2_1 _06633_ (.A(_02127_),
    .B(_02128_),
    .X(_02129_));
 sky130_fd_sc_hd__a21oi_1 _06634_ (.A1(_02109_),
    .A2(_02114_),
    .B1(_02129_),
    .Y(_02130_));
 sky130_fd_sc_hd__a31o_1 _06635_ (.A1(_02109_),
    .A2(_02114_),
    .A3(_02129_),
    .B1(_01789_),
    .X(_02131_));
 sky130_fd_sc_hd__a22o_1 _06636_ (.A1(\u_glbl_reg.reg_7[19] ),
    .A2(net610),
    .B1(net592),
    .B2(net169),
    .X(_02132_));
 sky130_fd_sc_hd__a211o_1 _06637_ (.A1(\u_glbl_reg.reg_23[19] ),
    .A2(net626),
    .B1(_01786_),
    .C1(_02132_),
    .X(_02133_));
 sky130_fd_sc_hd__a22o_1 _06638_ (.A1(\u_glbl_reg.reg_20[19] ),
    .A2(net640),
    .B1(net605),
    .B2(net209),
    .X(_02134_));
 sky130_fd_sc_hd__a221o_1 _06639_ (.A1(\u_glbl_reg.cfg_rst_ctrl[19] ),
    .A2(net701),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[19] ),
    .C1(_02134_),
    .X(_02135_));
 sky130_fd_sc_hd__a22o_1 _06640_ (.A1(\u_glbl_reg.reg_2[19] ),
    .A2(net687),
    .B1(net684),
    .B2(net475),
    .X(_02136_));
 sky130_fd_sc_hd__a221o_1 _06641_ (.A1(\u_glbl_reg.reg_17[19] ),
    .A2(net652),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[19] ),
    .C1(_02136_),
    .X(_02137_));
 sky130_fd_sc_hd__and3_1 _06642_ (.A(net1343),
    .B(\u_glbl_reg.reg_19[19] ),
    .C(net1139),
    .X(_02138_));
 sky130_fd_sc_hd__a221o_1 _06643_ (.A1(\u_glbl_reg.cfg_multi_func_sel[19] ),
    .A2(net618),
    .B1(net615),
    .B2(\u_glbl_reg.reg_6[19] ),
    .C1(_02138_),
    .X(_02139_));
 sky130_fd_sc_hd__a22o_1 _06644_ (.A1(\u_glbl_reg.reg_16[19] ),
    .A2(net1127),
    .B1(net635),
    .B2(\u_glbl_reg.reg_21[19] ),
    .X(_02140_));
 sky130_fd_sc_hd__a221o_1 _06645_ (.A1(\u_glbl_reg.reg_15[19] ),
    .A2(net658),
    .B1(net623),
    .B2(\u_glbl_reg.reg_3[19] ),
    .C1(_02140_),
    .X(_02141_));
 sky130_fd_sc_hd__or4_1 _06646_ (.A(_02135_),
    .B(_02137_),
    .C(_02139_),
    .D(_02141_),
    .X(_02142_));
 sky130_fd_sc_hd__a211oi_2 _06647_ (.A1(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ),
    .A2(net563),
    .B1(_02133_),
    .C1(_02142_),
    .Y(_02143_));
 sky130_fd_sc_hd__o21ai_1 _06648_ (.A1(net1985),
    .A2(_02131_),
    .B1(_02143_),
    .Y(\u_glbl_reg.reg_out[19] ));
 sky130_fd_sc_hd__or2_1 _06649_ (.A(net2122),
    .B(\u_glbl_reg.u_random.n0[20] ),
    .X(_02144_));
 sky130_fd_sc_hd__nand2_1 _06650_ (.A(net2122),
    .B(\u_glbl_reg.u_random.n0[20] ),
    .Y(_02145_));
 sky130_fd_sc_hd__and2_1 _06651_ (.A(_02144_),
    .B(_02145_),
    .X(_02146_));
 sky130_fd_sc_hd__or2_1 _06652_ (.A(_02110_),
    .B(_02129_),
    .X(_02147_));
 sky130_fd_sc_hd__o21ba_1 _06653_ (.A1(_02109_),
    .A2(_02128_),
    .B1_N(_02127_),
    .X(_02148_));
 sky130_fd_sc_hd__o21a_1 _06654_ (.A1(_02111_),
    .A2(_02147_),
    .B1(_02148_),
    .X(_02149_));
 sky130_fd_sc_hd__or2_1 _06655_ (.A(_02112_),
    .B(_02147_),
    .X(_02150_));
 sky130_fd_sc_hd__o21ai_2 _06656_ (.A1(_02074_),
    .A2(_02150_),
    .B1(_02149_),
    .Y(_02151_));
 sky130_fd_sc_hd__or2_1 _06657_ (.A(_02146_),
    .B(_02151_),
    .X(_02152_));
 sky130_fd_sc_hd__nand2_1 _06658_ (.A(_02146_),
    .B(_02151_),
    .Y(_02153_));
 sky130_fd_sc_hd__a22o_1 _06659_ (.A1(\u_glbl_reg.reg_19[20] ),
    .A2(net643),
    .B1(net631),
    .B2(\u_glbl_reg.reg_22[20] ),
    .X(_02154_));
 sky130_fd_sc_hd__a221o_1 _06660_ (.A1(\u_glbl_reg.reg_2[20] ),
    .A2(net689),
    .B1(net657),
    .B2(\u_glbl_reg.reg_15[20] ),
    .C1(_02154_),
    .X(_02155_));
 sky130_fd_sc_hd__a22o_1 _06661_ (.A1(\u_glbl_reg.reg_21[20] ),
    .A2(net635),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[20] ),
    .X(_02156_));
 sky130_fd_sc_hd__a211o_1 _06662_ (.A1(\u_glbl_reg.reg_20[20] ),
    .A2(net640),
    .B1(_02155_),
    .C1(_02156_),
    .X(_02157_));
 sky130_fd_sc_hd__a22o_1 _06663_ (.A1(\u_glbl_reg.reg_3[20] ),
    .A2(net623),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[20] ),
    .X(_02158_));
 sky130_fd_sc_hd__a221o_1 _06664_ (.A1(net477),
    .A2(net684),
    .B1(net562),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ),
    .C1(_02158_),
    .X(_02159_));
 sky130_fd_sc_hd__a22o_1 _06665_ (.A1(\u_glbl_reg.reg_23[20] ),
    .A2(net626),
    .B1(net592),
    .B2(net171),
    .X(_02160_));
 sky130_fd_sc_hd__a221o_1 _06666_ (.A1(\u_glbl_reg.cfg_rst_ctrl[20] ),
    .A2(net700),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[20] ),
    .C1(_02160_),
    .X(_02161_));
 sky130_fd_sc_hd__a22o_1 _06667_ (.A1(\u_glbl_reg.reg_16[20] ),
    .A2(net1127),
    .B1(net615),
    .B2(\u_glbl_reg.reg_6[20] ),
    .X(_02162_));
 sky130_fd_sc_hd__a221o_1 _06668_ (.A1(\u_glbl_reg.reg_17[20] ),
    .A2(net652),
    .B1(net605),
    .B2(net211),
    .C1(_02162_),
    .X(_02163_));
 sky130_fd_sc_hd__or4_1 _06669_ (.A(_02157_),
    .B(_02159_),
    .C(_02161_),
    .D(_02163_),
    .X(_02164_));
 sky130_fd_sc_hd__a31o_1 _06670_ (.A1(net593),
    .A2(_02152_),
    .A3(_02153_),
    .B1(_02164_),
    .X(\u_glbl_reg.reg_out[20] ));
 sky130_fd_sc_hd__and2_1 _06671_ (.A(\u_glbl_reg.u_random.n1_plus_n0[4] ),
    .B(\u_glbl_reg.u_random.n0[21] ),
    .X(_02165_));
 sky130_fd_sc_hd__nand2_1 _06672_ (.A(\u_glbl_reg.u_random.n1_plus_n0[4] ),
    .B(\u_glbl_reg.u_random.n0[21] ),
    .Y(_02166_));
 sky130_fd_sc_hd__nor2_1 _06673_ (.A(\u_glbl_reg.u_random.n1_plus_n0[4] ),
    .B(\u_glbl_reg.u_random.n0[21] ),
    .Y(_02167_));
 sky130_fd_sc_hd__or2_1 _06674_ (.A(_02165_),
    .B(_02167_),
    .X(_02168_));
 sky130_fd_sc_hd__a21bo_1 _06675_ (.A1(_02146_),
    .A2(_02151_),
    .B1_N(_02145_),
    .X(_02169_));
 sky130_fd_sc_hd__xnor2_1 _06676_ (.A(_02168_),
    .B(_02169_),
    .Y(_02170_));
 sky130_fd_sc_hd__a22o_1 _06677_ (.A1(\u_glbl_reg.reg_23[21] ),
    .A2(net626),
    .B1(net592),
    .B2(net172),
    .X(_02171_));
 sky130_fd_sc_hd__a221o_1 _06678_ (.A1(\u_glbl_reg.reg_19[21] ),
    .A2(net643),
    .B1(net605),
    .B2(net212),
    .C1(_02171_),
    .X(_02172_));
 sky130_fd_sc_hd__a22o_1 _06679_ (.A1(\u_glbl_reg.cfg_rst_ctrl[21] ),
    .A2(net701),
    .B1(net1127),
    .B2(\u_glbl_reg.reg_16[21] ),
    .X(_02173_));
 sky130_fd_sc_hd__a221o_1 _06680_ (.A1(\u_glbl_reg.reg_17[21] ),
    .A2(net653),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[21] ),
    .C1(_02173_),
    .X(_02174_));
 sky130_fd_sc_hd__a22o_1 _06681_ (.A1(net478),
    .A2(net684),
    .B1(net614),
    .B2(\u_glbl_reg.reg_6[21] ),
    .X(_02175_));
 sky130_fd_sc_hd__a221o_1 _06682_ (.A1(\u_glbl_reg.reg_2[21] ),
    .A2(net687),
    .B1(net648),
    .B2(\u_glbl_reg.reg_18[21] ),
    .C1(_02175_),
    .X(_02176_));
 sky130_fd_sc_hd__a22o_1 _06683_ (.A1(\u_glbl_reg.reg_21[21] ),
    .A2(net635),
    .B1(net619),
    .B2(\u_glbl_reg.cfg_multi_func_sel[21] ),
    .X(_02177_));
 sky130_fd_sc_hd__a22o_1 _06684_ (.A1(\u_glbl_reg.reg_15[21] ),
    .A2(net658),
    .B1(net631),
    .B2(\u_glbl_reg.reg_22[21] ),
    .X(_02178_));
 sky130_fd_sc_hd__a211o_1 _06685_ (.A1(\u_glbl_reg.reg_3[21] ),
    .A2(_01554_),
    .B1(_01786_),
    .C1(_02178_),
    .X(_02179_));
 sky130_fd_sc_hd__a211o_1 _06686_ (.A1(\u_glbl_reg.reg_20[21] ),
    .A2(net640),
    .B1(_02177_),
    .C1(_02179_),
    .X(_02180_));
 sky130_fd_sc_hd__a2111o_1 _06687_ (.A1(net2056),
    .A2(net562),
    .B1(_02174_),
    .C1(_02176_),
    .D1(_02180_),
    .X(_02181_));
 sky130_fd_sc_hd__a211o_1 _06688_ (.A1(net594),
    .A2(_02170_),
    .B1(_02172_),
    .C1(_02181_),
    .X(\u_glbl_reg.reg_out[21] ));
 sky130_fd_sc_hd__nand2_1 _06689_ (.A(net1995),
    .B(net1928),
    .Y(_02182_));
 sky130_fd_sc_hd__or2_1 _06690_ (.A(net1995),
    .B(\u_glbl_reg.u_random.n0[22] ),
    .X(_02183_));
 sky130_fd_sc_hd__nand2_1 _06691_ (.A(_02182_),
    .B(_02183_),
    .Y(_02184_));
 sky130_fd_sc_hd__a21o_1 _06692_ (.A1(_02145_),
    .A2(_02166_),
    .B1(_02167_),
    .X(_02185_));
 sky130_fd_sc_hd__nand4b_1 _06693_ (.A_N(_02168_),
    .B(_02151_),
    .C(_02145_),
    .D(_02144_),
    .Y(_02186_));
 sky130_fd_sc_hd__nand3_1 _06694_ (.A(_02184_),
    .B(_02185_),
    .C(_02186_),
    .Y(_02187_));
 sky130_fd_sc_hd__a21o_1 _06695_ (.A1(_02185_),
    .A2(_02186_),
    .B1(_02184_),
    .X(_02188_));
 sky130_fd_sc_hd__a22o_1 _06696_ (.A1(\u_glbl_reg.reg_16[22] ),
    .A2(net1127),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[22] ),
    .X(_02189_));
 sky130_fd_sc_hd__a22o_1 _06697_ (.A1(\u_glbl_reg.reg_23[22] ),
    .A2(net626),
    .B1(net623),
    .B2(\u_glbl_reg.reg_3[22] ),
    .X(_02190_));
 sky130_fd_sc_hd__a22o_1 _06698_ (.A1(\u_glbl_reg.reg_17[22] ),
    .A2(net652),
    .B1(net614),
    .B2(\u_glbl_reg.reg_6[22] ),
    .X(_02191_));
 sky130_fd_sc_hd__a221o_1 _06699_ (.A1(\u_glbl_reg.cfg_rst_ctrl[22] ),
    .A2(net701),
    .B1(net630),
    .B2(\u_glbl_reg.reg_22[22] ),
    .C1(_02190_),
    .X(_02192_));
 sky130_fd_sc_hd__a221o_1 _06700_ (.A1(\u_glbl_reg.reg_2[22] ),
    .A2(net689),
    .B1(net644),
    .B2(\u_glbl_reg.reg_19[22] ),
    .C1(_02189_),
    .X(_02193_));
 sky130_fd_sc_hd__a22o_1 _06701_ (.A1(net479),
    .A2(net684),
    .B1(net610),
    .B2(\u_glbl_reg.reg_7[22] ),
    .X(_02194_));
 sky130_fd_sc_hd__a221o_1 _06702_ (.A1(net213),
    .A2(net604),
    .B1(net591),
    .B2(net173),
    .C1(_02194_),
    .X(_02195_));
 sky130_fd_sc_hd__a211o_1 _06703_ (.A1(\u_glbl_reg.reg_15[22] ),
    .A2(net658),
    .B1(_01786_),
    .C1(_02191_),
    .X(_02196_));
 sky130_fd_sc_hd__a211o_1 _06704_ (.A1(\u_glbl_reg.reg_21[22] ),
    .A2(net635),
    .B1(_02195_),
    .C1(_02196_),
    .X(_02197_));
 sky130_fd_sc_hd__a221o_1 _06705_ (.A1(\u_glbl_reg.reg_20[22] ),
    .A2(net640),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[22] ),
    .C1(_02197_),
    .X(_02198_));
 sky130_fd_sc_hd__a211o_1 _06706_ (.A1(net2025),
    .A2(net562),
    .B1(_02193_),
    .C1(_02198_),
    .X(_02199_));
 sky130_fd_sc_hd__a311o_1 _06707_ (.A1(net593),
    .A2(_02187_),
    .A3(_02188_),
    .B1(_02192_),
    .C1(_02199_),
    .X(\u_glbl_reg.reg_out[22] ));
 sky130_fd_sc_hd__nor2_1 _06708_ (.A(\u_glbl_reg.u_random.n1_plus_n0[6] ),
    .B(\u_glbl_reg.u_random.n0[23] ),
    .Y(_02200_));
 sky130_fd_sc_hd__and2_1 _06709_ (.A(\u_glbl_reg.u_random.n1_plus_n0[6] ),
    .B(net1905),
    .X(_02201_));
 sky130_fd_sc_hd__or2_1 _06710_ (.A(_02200_),
    .B(_02201_),
    .X(_02202_));
 sky130_fd_sc_hd__a21oi_1 _06711_ (.A1(_02182_),
    .A2(_02188_),
    .B1(_02202_),
    .Y(_02203_));
 sky130_fd_sc_hd__a31o_1 _06712_ (.A1(_02182_),
    .A2(_02188_),
    .A3(_02202_),
    .B1(_01789_),
    .X(_02204_));
 sky130_fd_sc_hd__a22o_1 _06713_ (.A1(net480),
    .A2(net684),
    .B1(net626),
    .B2(\u_glbl_reg.reg_23[23] ),
    .X(_02205_));
 sky130_fd_sc_hd__a221o_1 _06714_ (.A1(\u_glbl_reg.cfg_rst_ctrl[23] ),
    .A2(net701),
    .B1(net562),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ),
    .C1(_02205_),
    .X(_02206_));
 sky130_fd_sc_hd__a22o_1 _06715_ (.A1(\u_glbl_reg.reg_20[23] ),
    .A2(net639),
    .B1(net618),
    .B2(\u_glbl_reg.cfg_multi_func_sel[23] ),
    .X(_02207_));
 sky130_fd_sc_hd__a22o_1 _06716_ (.A1(\u_glbl_reg.reg_19[23] ),
    .A2(net644),
    .B1(net605),
    .B2(net214),
    .X(_02208_));
 sky130_fd_sc_hd__a221o_1 _06717_ (.A1(\u_glbl_reg.reg_16[23] ),
    .A2(net1127),
    .B1(net615),
    .B2(\u_glbl_reg.reg_6[23] ),
    .C1(_02208_),
    .X(_02209_));
 sky130_fd_sc_hd__a2111o_1 _06718_ (.A1(\u_glbl_reg.reg_21[23] ),
    .A2(net635),
    .B1(_02206_),
    .C1(_02207_),
    .D1(_02209_),
    .X(_02210_));
 sky130_fd_sc_hd__a22o_1 _06719_ (.A1(\u_glbl_reg.reg_17[23] ),
    .A2(net653),
    .B1(net631),
    .B2(\u_glbl_reg.reg_22[23] ),
    .X(_02211_));
 sky130_fd_sc_hd__a221o_1 _06720_ (.A1(\u_glbl_reg.reg_3[23] ),
    .A2(net623),
    .B1(net611),
    .B2(\u_glbl_reg.reg_7[23] ),
    .C1(_02211_),
    .X(_02212_));
 sky130_fd_sc_hd__a22o_1 _06721_ (.A1(\u_glbl_reg.reg_15[23] ),
    .A2(net657),
    .B1(net647),
    .B2(\u_glbl_reg.reg_18[23] ),
    .X(_02213_));
 sky130_fd_sc_hd__a221o_1 _06722_ (.A1(\u_glbl_reg.reg_2[23] ),
    .A2(net687),
    .B1(net591),
    .B2(net174),
    .C1(_02213_),
    .X(_02214_));
 sky130_fd_sc_hd__nor3_1 _06723_ (.A(_02210_),
    .B(_02212_),
    .C(_02214_),
    .Y(_02215_));
 sky130_fd_sc_hd__o21ai_1 _06724_ (.A1(net1996),
    .A2(_02204_),
    .B1(_02215_),
    .Y(\u_glbl_reg.reg_out[23] ));
 sky130_fd_sc_hd__or2_1 _06725_ (.A(\u_glbl_reg.u_random.n1_plus_n0[7] ),
    .B(\u_glbl_reg.u_random.n0[24] ),
    .X(_02216_));
 sky130_fd_sc_hd__nand2_1 _06726_ (.A(\u_glbl_reg.u_random.n1_plus_n0[7] ),
    .B(net1892),
    .Y(_02217_));
 sky130_fd_sc_hd__and2_1 _06727_ (.A(_02216_),
    .B(_02217_),
    .X(_02218_));
 sky130_fd_sc_hd__or2_1 _06728_ (.A(_02184_),
    .B(_02202_),
    .X(_02219_));
 sky130_fd_sc_hd__or4b_2 _06729_ (.A(_02165_),
    .B(_02167_),
    .C(_02219_),
    .D_N(_02146_),
    .X(_02220_));
 sky130_fd_sc_hd__o21ba_1 _06730_ (.A1(_02182_),
    .A2(_02200_),
    .B1_N(_02201_),
    .X(_02221_));
 sky130_fd_sc_hd__o221a_1 _06731_ (.A1(_02185_),
    .A2(_02219_),
    .B1(_02220_),
    .B2(_02149_),
    .C1(_02221_),
    .X(_02222_));
 sky130_fd_sc_hd__o31ai_4 _06732_ (.A1(_02074_),
    .A2(_02150_),
    .A3(_02220_),
    .B1(_02222_),
    .Y(_02223_));
 sky130_fd_sc_hd__nand2_1 _06733_ (.A(_02218_),
    .B(_02223_),
    .Y(_02224_));
 sky130_fd_sc_hd__o21a_1 _06734_ (.A1(_02218_),
    .A2(_02223_),
    .B1(net593),
    .X(_02225_));
 sky130_fd_sc_hd__a22o_1 _06735_ (.A1(\u_glbl_reg.reg_2[24] ),
    .A2(net685),
    .B1(net633),
    .B2(\u_glbl_reg.reg_21[24] ),
    .X(_02226_));
 sky130_fd_sc_hd__a221o_1 _06736_ (.A1(\u_glbl_reg.cfg_rst_ctrl[24] ),
    .A2(net699),
    .B1(net641),
    .B2(\u_glbl_reg.reg_19[24] ),
    .C1(_02226_),
    .X(_02227_));
 sky130_fd_sc_hd__a22o_1 _06737_ (.A1(\u_glbl_reg.reg_3[24] ),
    .A2(net620),
    .B1(net607),
    .B2(\u_glbl_reg.reg_7[24] ),
    .X(_02228_));
 sky130_fd_sc_hd__a22o_1 _06738_ (.A1(\u_glbl_reg.reg_15[24] ),
    .A2(net654),
    .B1(net589),
    .B2(net175),
    .X(_02229_));
 sky130_fd_sc_hd__a22o_1 _06739_ (.A1(net481),
    .A2(net681),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[24] ),
    .X(_02230_));
 sky130_fd_sc_hd__a22o_1 _06740_ (.A1(\u_glbl_reg.reg_18[24] ),
    .A2(net645),
    .B1(net616),
    .B2(\u_glbl_reg.cfg_multi_func_sel[24] ),
    .X(_02231_));
 sky130_fd_sc_hd__a221o_1 _06741_ (.A1(\u_glbl_reg.reg_16[24] ),
    .A2(net1124),
    .B1(net624),
    .B2(\u_glbl_reg.reg_23[24] ),
    .C1(_02231_),
    .X(_02232_));
 sky130_fd_sc_hd__a22o_1 _06742_ (.A1(\u_glbl_reg.reg_20[24] ),
    .A2(net637),
    .B1(net603),
    .B2(net1107),
    .X(_02233_));
 sky130_fd_sc_hd__a221o_1 _06743_ (.A1(\u_glbl_reg.reg_17[24] ),
    .A2(net649),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[24] ),
    .C1(_02233_),
    .X(_02234_));
 sky130_fd_sc_hd__or4_1 _06744_ (.A(_02229_),
    .B(_02230_),
    .C(_02232_),
    .D(_02234_),
    .X(_02235_));
 sky130_fd_sc_hd__a2111o_2 _06745_ (.A1(net2014),
    .A2(net560),
    .B1(_02227_),
    .C1(_02228_),
    .D1(_02235_),
    .X(_02236_));
 sky130_fd_sc_hd__a21o_1 _06746_ (.A1(_02224_),
    .A2(_02225_),
    .B1(_02236_),
    .X(\u_glbl_reg.reg_out[24] ));
 sky130_fd_sc_hd__nor2_1 _06747_ (.A(\u_glbl_reg.u_random.n1_plus_n0[8] ),
    .B(\u_glbl_reg.u_random.n0[25] ),
    .Y(_02237_));
 sky130_fd_sc_hd__nand2_1 _06748_ (.A(\u_glbl_reg.u_random.n1_plus_n0[8] ),
    .B(\u_glbl_reg.u_random.n0[25] ),
    .Y(_02238_));
 sky130_fd_sc_hd__and2b_1 _06749_ (.A_N(_02237_),
    .B(_02238_),
    .X(_02239_));
 sky130_fd_sc_hd__a21bo_1 _06750_ (.A1(_02218_),
    .A2(_02223_),
    .B1_N(_02217_),
    .X(_02240_));
 sky130_fd_sc_hd__xnor2_1 _06751_ (.A(_02239_),
    .B(_02240_),
    .Y(_02241_));
 sky130_fd_sc_hd__nor2_2 _06752_ (.A(_01789_),
    .B(_02241_),
    .Y(_02242_));
 sky130_fd_sc_hd__a22o_1 _06753_ (.A1(net482),
    .A2(net681),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[25] ),
    .X(_02243_));
 sky130_fd_sc_hd__a221o_1 _06754_ (.A1(\u_glbl_reg.reg_2[25] ),
    .A2(net685),
    .B1(net560),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ),
    .C1(_02243_),
    .X(_02244_));
 sky130_fd_sc_hd__a22o_1 _06755_ (.A1(\u_glbl_reg.reg_20[25] ),
    .A2(net637),
    .B1(net633),
    .B2(\u_glbl_reg.reg_21[25] ),
    .X(_02245_));
 sky130_fd_sc_hd__a22o_1 _06756_ (.A1(\u_glbl_reg.reg_15[25] ),
    .A2(net654),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[25] ),
    .X(_02246_));
 sky130_fd_sc_hd__a211o_1 _06757_ (.A1(\u_glbl_reg.reg_3[25] ),
    .A2(net620),
    .B1(_01786_),
    .C1(_02246_),
    .X(_02247_));
 sky130_fd_sc_hd__a2111o_1 _06758_ (.A1(\u_glbl_reg.cfg_multi_func_sel[25] ),
    .A2(net616),
    .B1(_02244_),
    .C1(_02245_),
    .D1(_02247_),
    .X(_02248_));
 sky130_fd_sc_hd__a22o_1 _06759_ (.A1(\u_glbl_reg.reg_23[25] ),
    .A2(net624),
    .B1(net589),
    .B2(net176),
    .X(_02249_));
 sky130_fd_sc_hd__a221o_1 _06760_ (.A1(\u_glbl_reg.reg_19[25] ),
    .A2(net641),
    .B1(net603),
    .B2(net1106),
    .C1(_02249_),
    .X(_02250_));
 sky130_fd_sc_hd__a22o_1 _06761_ (.A1(\u_glbl_reg.cfg_rst_ctrl[25] ),
    .A2(net699),
    .B1(net1124),
    .B2(\u_glbl_reg.reg_16[25] ),
    .X(_02251_));
 sky130_fd_sc_hd__a22o_1 _06762_ (.A1(\u_glbl_reg.reg_18[25] ),
    .A2(net646),
    .B1(net607),
    .B2(\u_glbl_reg.reg_7[25] ),
    .X(_02252_));
 sky130_fd_sc_hd__a2111o_1 _06763_ (.A1(net2278),
    .A2(net649),
    .B1(_02250_),
    .C1(_02251_),
    .D1(_02252_),
    .X(_02253_));
 sky130_fd_sc_hd__or3_1 _06764_ (.A(_02242_),
    .B(_02248_),
    .C(_02253_),
    .X(\u_glbl_reg.reg_out[25] ));
 sky130_fd_sc_hd__or2_1 _06765_ (.A(net2003),
    .B(net1915),
    .X(_02254_));
 sky130_fd_sc_hd__nand2_1 _06766_ (.A(net2003),
    .B(net1915),
    .Y(_02255_));
 sky130_fd_sc_hd__and3_1 _06767_ (.A(_02218_),
    .B(_02223_),
    .C(_02239_),
    .X(_02256_));
 sky130_fd_sc_hd__a21oi_1 _06768_ (.A1(_02217_),
    .A2(_02238_),
    .B1(_02237_),
    .Y(_02257_));
 sky130_fd_sc_hd__a211o_1 _06769_ (.A1(_02254_),
    .A2(_02255_),
    .B1(_02256_),
    .C1(_02257_),
    .X(_02258_));
 sky130_fd_sc_hd__o211ai_2 _06770_ (.A1(_02256_),
    .A2(_02257_),
    .B1(_02254_),
    .C1(_02255_),
    .Y(_02259_));
 sky130_fd_sc_hd__a22o_1 _06771_ (.A1(\u_glbl_reg.reg_16[26] ),
    .A2(net1126),
    .B1(net651),
    .B2(\u_glbl_reg.reg_17[26] ),
    .X(_02260_));
 sky130_fd_sc_hd__a22o_1 _06772_ (.A1(\u_glbl_reg.reg_19[26] ),
    .A2(net642),
    .B1(net632),
    .B2(\u_glbl_reg.reg_22[26] ),
    .X(_02261_));
 sky130_fd_sc_hd__a22o_1 _06773_ (.A1(net483),
    .A2(net681),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[26] ),
    .X(_02262_));
 sky130_fd_sc_hd__a221o_1 _06774_ (.A1(\u_glbl_reg.reg_23[26] ),
    .A2(net624),
    .B1(net589),
    .B2(net177),
    .C1(_02262_),
    .X(_02263_));
 sky130_fd_sc_hd__a22o_1 _06775_ (.A1(\u_glbl_reg.reg_3[26] ),
    .A2(net620),
    .B1(net604),
    .B2(net1105),
    .X(_02264_));
 sky130_fd_sc_hd__a221o_1 _06776_ (.A1(\u_glbl_reg.reg_7[26] ),
    .A2(net607),
    .B1(net560),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ),
    .C1(_02264_),
    .X(_02265_));
 sky130_fd_sc_hd__a22o_1 _06777_ (.A1(\u_glbl_reg.cfg_rst_ctrl[26] ),
    .A2(net698),
    .B1(net645),
    .B2(\u_glbl_reg.reg_18[26] ),
    .X(_02266_));
 sky130_fd_sc_hd__a221o_1 _06778_ (.A1(\u_glbl_reg.reg_2[26] ),
    .A2(net685),
    .B1(net654),
    .B2(\u_glbl_reg.reg_15[26] ),
    .C1(_02266_),
    .X(_02267_));
 sky130_fd_sc_hd__a22o_1 _06779_ (.A1(\u_glbl_reg.reg_20[26] ),
    .A2(net637),
    .B1(net616),
    .B2(\u_glbl_reg.cfg_multi_func_sel[26] ),
    .X(_02268_));
 sky130_fd_sc_hd__a21o_1 _06780_ (.A1(\u_glbl_reg.reg_21[26] ),
    .A2(net633),
    .B1(_02268_),
    .X(_02269_));
 sky130_fd_sc_hd__or4_2 _06781_ (.A(_02263_),
    .B(_02265_),
    .C(_02267_),
    .D(_02269_),
    .X(_02270_));
 sky130_fd_sc_hd__or3_4 _06782_ (.A(_02260_),
    .B(_02261_),
    .C(_02270_),
    .X(_02271_));
 sky130_fd_sc_hd__a31o_1 _06783_ (.A1(net593),
    .A2(_02258_),
    .A3(net2004),
    .B1(_02271_),
    .X(\u_glbl_reg.reg_out[26] ));
 sky130_fd_sc_hd__nor2_1 _06784_ (.A(net2036),
    .B(net1894),
    .Y(_02272_));
 sky130_fd_sc_hd__and2_1 _06785_ (.A(net2036),
    .B(net1894),
    .X(_02273_));
 sky130_fd_sc_hd__a211o_1 _06786_ (.A1(_02255_),
    .A2(_02259_),
    .B1(_02272_),
    .C1(_02273_),
    .X(_02274_));
 sky130_fd_sc_hd__o211ai_1 _06787_ (.A1(_02272_),
    .A2(_02273_),
    .B1(_02255_),
    .C1(_02259_),
    .Y(_02275_));
 sky130_fd_sc_hd__a22o_1 _06788_ (.A1(\u_glbl_reg.cfg_rst_ctrl[27] ),
    .A2(net698),
    .B1(net645),
    .B2(\u_glbl_reg.reg_18[27] ),
    .X(_02276_));
 sky130_fd_sc_hd__a22o_1 _06789_ (.A1(\u_glbl_reg.reg_20[27] ),
    .A2(net637),
    .B1(net616),
    .B2(\u_glbl_reg.cfg_multi_func_sel[27] ),
    .X(_02277_));
 sky130_fd_sc_hd__a22o_1 _06790_ (.A1(\u_glbl_reg.reg_19[27] ),
    .A2(net641),
    .B1(net604),
    .B2(net1104),
    .X(_02278_));
 sky130_fd_sc_hd__a221o_1 _06791_ (.A1(\u_glbl_reg.reg_16[27] ),
    .A2(net1124),
    .B1(net613),
    .B2(\u_glbl_reg.reg_6[27] ),
    .C1(_02278_),
    .X(_02279_));
 sky130_fd_sc_hd__a211o_1 _06792_ (.A1(\u_glbl_reg.reg_21[27] ),
    .A2(net633),
    .B1(_02277_),
    .C1(_02279_),
    .X(_02280_));
 sky130_fd_sc_hd__a22o_1 _06793_ (.A1(net484),
    .A2(net681),
    .B1(net624),
    .B2(\u_glbl_reg.reg_23[27] ),
    .X(_02281_));
 sky130_fd_sc_hd__a221o_1 _06794_ (.A1(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ),
    .A2(net560),
    .B1(net589),
    .B2(net178),
    .C1(_02281_),
    .X(_02282_));
 sky130_fd_sc_hd__a221o_1 _06795_ (.A1(\u_glbl_reg.reg_2[27] ),
    .A2(net685),
    .B1(net654),
    .B2(\u_glbl_reg.reg_15[27] ),
    .C1(_02276_),
    .X(_02283_));
 sky130_fd_sc_hd__a22o_1 _06796_ (.A1(\u_glbl_reg.reg_17[27] ),
    .A2(net649),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[27] ),
    .X(_02284_));
 sky130_fd_sc_hd__a221o_1 _06797_ (.A1(\u_glbl_reg.reg_3[27] ),
    .A2(net620),
    .B1(net607),
    .B2(\u_glbl_reg.reg_7[27] ),
    .C1(_02284_),
    .X(_02285_));
 sky130_fd_sc_hd__or4_4 _06798_ (.A(_02280_),
    .B(_02282_),
    .C(_02283_),
    .D(_02285_),
    .X(_02286_));
 sky130_fd_sc_hd__a31o_1 _06799_ (.A1(net593),
    .A2(_02274_),
    .A3(_02275_),
    .B1(_02286_),
    .X(\u_glbl_reg.reg_out[27] ));
 sky130_fd_sc_hd__xnor2_1 _06800_ (.A(net2018),
    .B(net1897),
    .Y(_02287_));
 sky130_fd_sc_hd__nor2_1 _06801_ (.A(_02255_),
    .B(_02272_),
    .Y(_02288_));
 sky130_fd_sc_hd__or3_1 _06802_ (.A(_02257_),
    .B(_02273_),
    .C(_02288_),
    .X(_02289_));
 sky130_fd_sc_hd__a31o_1 _06803_ (.A1(_02218_),
    .A2(_02223_),
    .A3(_02239_),
    .B1(_02289_),
    .X(_02290_));
 sky130_fd_sc_hd__o21ba_1 _06804_ (.A1(_02254_),
    .A2(_02273_),
    .B1_N(_02272_),
    .X(_02291_));
 sky130_fd_sc_hd__a21bo_1 _06805_ (.A1(_02290_),
    .A2(_02291_),
    .B1_N(_02287_),
    .X(_02292_));
 sky130_fd_sc_hd__and3b_1 _06806_ (.A_N(_02287_),
    .B(_02290_),
    .C(_02291_),
    .X(_02293_));
 sky130_fd_sc_hd__nor2_1 _06807_ (.A(_01789_),
    .B(_02293_),
    .Y(_02294_));
 sky130_fd_sc_hd__a22o_1 _06808_ (.A1(\u_glbl_reg.reg_19[28] ),
    .A2(net641),
    .B1(net624),
    .B2(\u_glbl_reg.reg_23[28] ),
    .X(_02295_));
 sky130_fd_sc_hd__a22o_1 _06809_ (.A1(\u_glbl_reg.reg_17[28] ),
    .A2(net649),
    .B1(net645),
    .B2(\u_glbl_reg.reg_18[28] ),
    .X(_02296_));
 sky130_fd_sc_hd__a221o_1 _06810_ (.A1(\u_glbl_reg.reg_15[28] ),
    .A2(net654),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[28] ),
    .C1(_02296_),
    .X(_02297_));
 sky130_fd_sc_hd__a22o_1 _06811_ (.A1(\u_glbl_reg.reg_20[28] ),
    .A2(net637),
    .B1(net616),
    .B2(\u_glbl_reg.cfg_multi_func_sel[28] ),
    .X(_02298_));
 sky130_fd_sc_hd__a211o_1 _06812_ (.A1(\u_glbl_reg.reg_21[28] ),
    .A2(net633),
    .B1(_02297_),
    .C1(_02298_),
    .X(_02299_));
 sky130_fd_sc_hd__a22o_1 _06813_ (.A1(net485),
    .A2(net681),
    .B1(net1124),
    .B2(\u_glbl_reg.reg_16[28] ),
    .X(_02300_));
 sky130_fd_sc_hd__a221o_1 _06814_ (.A1(\u_glbl_reg.reg_7[28] ),
    .A2(net607),
    .B1(net560),
    .B2(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ),
    .C1(_02300_),
    .X(_02301_));
 sky130_fd_sc_hd__a22o_1 _06815_ (.A1(\u_glbl_reg.reg_2[28] ),
    .A2(net685),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[28] ),
    .X(_02302_));
 sky130_fd_sc_hd__a221o_1 _06816_ (.A1(\u_glbl_reg.cfg_rst_ctrl[28] ),
    .A2(net698),
    .B1(net603),
    .B2(net1103),
    .C1(_02302_),
    .X(_02303_));
 sky130_fd_sc_hd__a221o_1 _06817_ (.A1(\u_glbl_reg.reg_3[28] ),
    .A2(net620),
    .B1(net590),
    .B2(net179),
    .C1(_02295_),
    .X(_02304_));
 sky130_fd_sc_hd__or4_4 _06818_ (.A(_02299_),
    .B(_02301_),
    .C(_02303_),
    .D(_02304_),
    .X(_02305_));
 sky130_fd_sc_hd__a21o_1 _06819_ (.A1(net2019),
    .A2(_02294_),
    .B1(_02305_),
    .X(\u_glbl_reg.reg_out[28] ));
 sky130_fd_sc_hd__or2_1 _06820_ (.A(\u_glbl_reg.u_random.n1_plus_n0[12] ),
    .B(\u_glbl_reg.u_random.n0[29] ),
    .X(_02306_));
 sky130_fd_sc_hd__nand2_1 _06821_ (.A(\u_glbl_reg.u_random.n1_plus_n0[12] ),
    .B(\u_glbl_reg.u_random.n0[29] ),
    .Y(_02307_));
 sky130_fd_sc_hd__nand2_2 _06822_ (.A(_02306_),
    .B(_02307_),
    .Y(_02308_));
 sky130_fd_sc_hd__a21o_1 _06823_ (.A1(\u_glbl_reg.u_random.n1_plus_n0[11] ),
    .A2(\u_glbl_reg.u_random.n0[28] ),
    .B1(_02293_),
    .X(_02309_));
 sky130_fd_sc_hd__xnor2_4 _06824_ (.A(_02308_),
    .B(_02309_),
    .Y(_02310_));
 sky130_fd_sc_hd__a22o_1 _06825_ (.A1(\u_glbl_reg.reg_17[29] ),
    .A2(net651),
    .B1(net629),
    .B2(\u_glbl_reg.reg_22[29] ),
    .X(_02311_));
 sky130_fd_sc_hd__a22o_1 _06826_ (.A1(\u_glbl_reg.reg_19[29] ),
    .A2(net642),
    .B1(net603),
    .B2(net1102),
    .X(_02312_));
 sky130_fd_sc_hd__a22o_1 _06827_ (.A1(\u_glbl_reg.cfg_rst_ctrl[29] ),
    .A2(net698),
    .B1(net685),
    .B2(\u_glbl_reg.reg_2[29] ),
    .X(_02313_));
 sky130_fd_sc_hd__a221o_1 _06828_ (.A1(\u_glbl_reg.reg_15[29] ),
    .A2(net654),
    .B1(net645),
    .B2(\u_glbl_reg.reg_18[29] ),
    .C1(_02313_),
    .X(_02314_));
 sky130_fd_sc_hd__a221o_1 _06829_ (.A1(\u_glbl_reg.reg_3[29] ),
    .A2(net620),
    .B1(net609),
    .B2(\u_glbl_reg.reg_7[29] ),
    .C1(_02312_),
    .X(_02315_));
 sky130_fd_sc_hd__a22o_1 _06830_ (.A1(net486),
    .A2(net681),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[29] ),
    .X(_02316_));
 sky130_fd_sc_hd__a221o_1 _06831_ (.A1(\u_glbl_reg.reg_23[29] ),
    .A2(net624),
    .B1(net589),
    .B2(net180),
    .C1(_02316_),
    .X(_02317_));
 sky130_fd_sc_hd__a211o_1 _06832_ (.A1(\u_glbl_reg.cfg_multi_func_sel[29] ),
    .A2(net616),
    .B1(_02314_),
    .C1(_02317_),
    .X(_02318_));
 sky130_fd_sc_hd__a221o_1 _06833_ (.A1(\u_glbl_reg.reg_20[29] ),
    .A2(net637),
    .B1(net633),
    .B2(\u_glbl_reg.reg_21[29] ),
    .C1(_02318_),
    .X(_02319_));
 sky130_fd_sc_hd__a221o_1 _06834_ (.A1(net2001),
    .A2(net560),
    .B1(net595),
    .B2(_02310_),
    .C1(_02319_),
    .X(_02320_));
 sky130_fd_sc_hd__a2111o_1 _06835_ (.A1(\u_glbl_reg.reg_16[29] ),
    .A2(net1126),
    .B1(_02311_),
    .C1(_02315_),
    .D1(_02320_),
    .X(\u_glbl_reg.reg_out[29] ));
 sky130_fd_sc_hd__and2_1 _06836_ (.A(\u_glbl_reg.u_random.n1_plus_n0[13] ),
    .B(\u_glbl_reg.u_random.n0[30] ),
    .X(_02321_));
 sky130_fd_sc_hd__nor2_1 _06837_ (.A(\u_glbl_reg.u_random.n1_plus_n0[13] ),
    .B(\u_glbl_reg.u_random.n0[30] ),
    .Y(_02322_));
 sky130_fd_sc_hd__nor2_1 _06838_ (.A(_02321_),
    .B(_02322_),
    .Y(_02323_));
 sky130_fd_sc_hd__a22o_1 _06839_ (.A1(\u_glbl_reg.u_random.n1_plus_n0[11] ),
    .A2(\u_glbl_reg.u_random.n0[28] ),
    .B1(\u_glbl_reg.u_random.n1_plus_n0[12] ),
    .B2(\u_glbl_reg.u_random.n0[29] ),
    .X(_02324_));
 sky130_fd_sc_hd__o21a_1 _06840_ (.A1(_02293_),
    .A2(_02324_),
    .B1(_02306_),
    .X(_02325_));
 sky130_fd_sc_hd__xnor2_2 _06841_ (.A(_02323_),
    .B(_02325_),
    .Y(_02326_));
 sky130_fd_sc_hd__nor2_4 _06842_ (.A(_01789_),
    .B(_02326_),
    .Y(_02327_));
 sky130_fd_sc_hd__a22o_1 _06843_ (.A1(\u_glbl_reg.reg_23[30] ),
    .A2(net624),
    .B1(net612),
    .B2(\u_glbl_reg.reg_6[30] ),
    .X(_02328_));
 sky130_fd_sc_hd__a221o_1 _06844_ (.A1(\u_glbl_reg.reg_15[30] ),
    .A2(net654),
    .B1(net637),
    .B2(\u_glbl_reg.reg_20[30] ),
    .C1(_02328_),
    .X(_02329_));
 sky130_fd_sc_hd__a22o_1 _06845_ (.A1(\u_glbl_reg.reg_2[30] ),
    .A2(net685),
    .B1(net1124),
    .B2(\u_glbl_reg.reg_16[30] ),
    .X(_02330_));
 sky130_fd_sc_hd__a211o_1 _06846_ (.A1(net2035),
    .A2(net560),
    .B1(_02329_),
    .C1(_02330_),
    .X(_02331_));
 sky130_fd_sc_hd__a22o_1 _06847_ (.A1(\u_glbl_reg.reg_21[30] ),
    .A2(net633),
    .B1(net620),
    .B2(\u_glbl_reg.reg_3[30] ),
    .X(_02332_));
 sky130_fd_sc_hd__a221o_1 _06848_ (.A1(\u_glbl_reg.reg_22[30] ),
    .A2(net628),
    .B1(net607),
    .B2(\u_glbl_reg.reg_7[30] ),
    .C1(_02332_),
    .X(_02333_));
 sky130_fd_sc_hd__a22o_1 _06849_ (.A1(\u_glbl_reg.reg_19[30] ),
    .A2(net644),
    .B1(net603),
    .B2(net1101),
    .X(_02334_));
 sky130_fd_sc_hd__a221o_1 _06850_ (.A1(\u_glbl_reg.cfg_rst_ctrl[30] ),
    .A2(net699),
    .B1(net683),
    .B2(net488),
    .C1(_02334_),
    .X(_02335_));
 sky130_fd_sc_hd__a22o_1 _06851_ (.A1(\u_glbl_reg.reg_17[30] ),
    .A2(net649),
    .B1(net590),
    .B2(net182),
    .X(_02336_));
 sky130_fd_sc_hd__a221o_1 _06852_ (.A1(\u_glbl_reg.reg_18[30] ),
    .A2(net646),
    .B1(net616),
    .B2(net1109),
    .C1(_02336_),
    .X(_02337_));
 sky130_fd_sc_hd__or3_1 _06853_ (.A(_02333_),
    .B(_02335_),
    .C(_02337_),
    .X(_02338_));
 sky130_fd_sc_hd__or3_2 _06854_ (.A(_02327_),
    .B(_02331_),
    .C(_02338_),
    .X(\u_glbl_reg.reg_out[30] ));
 sky130_fd_sc_hd__a21o_1 _06855_ (.A1(_02323_),
    .A2(_02325_),
    .B1(_02321_),
    .X(_02339_));
 sky130_fd_sc_hd__xnor2_2 _06856_ (.A(\u_glbl_reg.u_random.n1_plus_n0[14] ),
    .B(\u_glbl_reg.u_random.n0[31] ),
    .Y(_02340_));
 sky130_fd_sc_hd__xnor2_4 _06857_ (.A(_02339_),
    .B(_02340_),
    .Y(_02341_));
 sky130_fd_sc_hd__a22o_1 _06858_ (.A1(\u_glbl_reg.reg_3[31] ),
    .A2(net620),
    .B1(net609),
    .B2(\u_glbl_reg.reg_7[31] ),
    .X(_02342_));
 sky130_fd_sc_hd__a22o_1 _06859_ (.A1(\u_glbl_reg.reg_19[31] ),
    .A2(net641),
    .B1(_01553_),
    .B2(\u_glbl_reg.reg_23[31] ),
    .X(_02343_));
 sky130_fd_sc_hd__a221o_1 _06860_ (.A1(\u_glbl_reg.reg_16[31] ),
    .A2(net1124),
    .B1(net615),
    .B2(\u_glbl_reg.reg_6[31] ),
    .C1(_02342_),
    .X(_02344_));
 sky130_fd_sc_hd__a22o_1 _06861_ (.A1(net489),
    .A2(net681),
    .B1(net628),
    .B2(\u_glbl_reg.reg_22[31] ),
    .X(_02345_));
 sky130_fd_sc_hd__a221o_1 _06862_ (.A1(\u_glbl_reg.reg_2[31] ),
    .A2(net685),
    .B1(net654),
    .B2(\u_glbl_reg.reg_15[31] ),
    .C1(_02345_),
    .X(_02346_));
 sky130_fd_sc_hd__a22o_1 _06863_ (.A1(net1100),
    .A2(net603),
    .B1(net590),
    .B2(net183),
    .X(_02347_));
 sky130_fd_sc_hd__a221o_1 _06864_ (.A1(\u_glbl_reg.reg_17[31] ),
    .A2(net649),
    .B1(net646),
    .B2(\u_glbl_reg.reg_18[31] ),
    .C1(_02347_),
    .X(_02348_));
 sky130_fd_sc_hd__a211o_1 _06865_ (.A1(\u_glbl_reg.cfg_rst_ctrl[31] ),
    .A2(net699),
    .B1(_01786_),
    .C1(_02343_),
    .X(_02349_));
 sky130_fd_sc_hd__a211o_1 _06866_ (.A1(\u_glbl_reg.reg_20[31] ),
    .A2(net637),
    .B1(_02348_),
    .C1(_02349_),
    .X(_02350_));
 sky130_fd_sc_hd__a221o_1 _06867_ (.A1(\u_glbl_reg.reg_21[31] ),
    .A2(net633),
    .B1(net616),
    .B2(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .C1(_02350_),
    .X(_02351_));
 sky130_fd_sc_hd__a211o_1 _06868_ (.A1(net2065),
    .A2(net560),
    .B1(_02346_),
    .C1(_02351_),
    .X(_02352_));
 sky130_fd_sc_hd__a211o_1 _06869_ (.A1(net595),
    .A2(_02341_),
    .B1(_02344_),
    .C1(_02352_),
    .X(\u_glbl_reg.reg_out[31] ));
 sky130_fd_sc_hd__and3_1 _06870_ (.A(net1360),
    .B(net1261),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[0] ),
    .X(_02353_));
 sky130_fd_sc_hd__a221o_1 _06871_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[0] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[0] ),
    .C1(net1246),
    .X(_02354_));
 sky130_fd_sc_hd__o22a_1 _06872_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[0] ),
    .A2(net1230),
    .B1(_02353_),
    .B2(_02354_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__and3_1 _06873_ (.A(net1360),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ),
    .X(_02355_));
 sky130_fd_sc_hd__a221o_1 _06874_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[1] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[1] ),
    .C1(net1246),
    .X(_02356_));
 sky130_fd_sc_hd__o22a_1 _06875_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[1] ),
    .A2(net1230),
    .B1(_02355_),
    .B2(_02356_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__and3_1 _06876_ (.A(net1360),
    .B(net1261),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[2] ),
    .X(_02357_));
 sky130_fd_sc_hd__a221o_1 _06877_ (.A1(net1285),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[2] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ),
    .C1(net1246),
    .X(_02358_));
 sky130_fd_sc_hd__o22a_1 _06878_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[2] ),
    .A2(net1230),
    .B1(_02357_),
    .B2(_02358_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__and3_1 _06879_ (.A(net1360),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ),
    .X(_02359_));
 sky130_fd_sc_hd__a221o_1 _06880_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[3] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[3] ),
    .C1(net1246),
    .X(_02360_));
 sky130_fd_sc_hd__o22a_1 _06881_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[3] ),
    .A2(net1230),
    .B1(_02359_),
    .B2(_02360_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__and3_1 _06882_ (.A(net1360),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ),
    .X(_02361_));
 sky130_fd_sc_hd__a221o_1 _06883_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[4] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[4] ),
    .C1(net1243),
    .X(_02362_));
 sky130_fd_sc_hd__o22a_1 _06884_ (.A1(net2166),
    .A2(net1230),
    .B1(_02361_),
    .B2(_02362_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__and3_1 _06885_ (.A(net1360),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ),
    .X(_02363_));
 sky130_fd_sc_hd__a221o_1 _06886_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[5] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[5] ),
    .C1(net1243),
    .X(_02364_));
 sky130_fd_sc_hd__o22a_1 _06887_ (.A1(net2266),
    .A2(net1230),
    .B1(_02363_),
    .B2(_02364_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__and3_1 _06888_ (.A(net1361),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ),
    .X(_02365_));
 sky130_fd_sc_hd__a221o_1 _06889_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[6] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[6] ),
    .C1(net1243),
    .X(_02366_));
 sky130_fd_sc_hd__o22a_1 _06890_ (.A1(net2349),
    .A2(net1230),
    .B1(_02365_),
    .B2(_02366_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__and3_1 _06891_ (.A(net1354),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ),
    .X(_02367_));
 sky130_fd_sc_hd__a221o_1 _06892_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[7] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[7] ),
    .C1(net1246),
    .X(_02368_));
 sky130_fd_sc_hd__o22a_1 _06893_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[7] ),
    .A2(net1229),
    .B1(_02367_),
    .B2(_02368_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__and3_1 _06894_ (.A(net1354),
    .B(net1260),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[8] ),
    .X(_02369_));
 sky130_fd_sc_hd__a221o_1 _06895_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[8] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ),
    .C1(net1245),
    .X(_02370_));
 sky130_fd_sc_hd__o22a_1 _06896_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[8] ),
    .A2(net1229),
    .B1(_02369_),
    .B2(_02370_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__and3_1 _06897_ (.A(net1354),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ),
    .X(_02371_));
 sky130_fd_sc_hd__a221o_1 _06898_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[9] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[9] ),
    .C1(net1244),
    .X(_02372_));
 sky130_fd_sc_hd__o22a_1 _06899_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[9] ),
    .A2(net1229),
    .B1(_02371_),
    .B2(_02372_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__and3_1 _06900_ (.A(net1354),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ),
    .X(_02373_));
 sky130_fd_sc_hd__a221o_1 _06901_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[10] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[10] ),
    .C1(net1244),
    .X(_02374_));
 sky130_fd_sc_hd__o22a_1 _06902_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[10] ),
    .A2(net1229),
    .B1(_02373_),
    .B2(_02374_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__and3_1 _06903_ (.A(net1354),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ),
    .X(_02375_));
 sky130_fd_sc_hd__a221o_1 _06904_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[11] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[11] ),
    .C1(net1244),
    .X(_02376_));
 sky130_fd_sc_hd__o22a_1 _06905_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[11] ),
    .A2(net1229),
    .B1(_02375_),
    .B2(_02376_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__and3_1 _06906_ (.A(net1354),
    .B(net1260),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[12] ),
    .X(_02377_));
 sky130_fd_sc_hd__a221o_1 _06907_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[12] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ),
    .C1(net1243),
    .X(_02378_));
 sky130_fd_sc_hd__o22a_1 _06908_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[12] ),
    .A2(net1229),
    .B1(_02377_),
    .B2(_02378_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__and3_1 _06909_ (.A(net1354),
    .B(net1367),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ),
    .X(_02379_));
 sky130_fd_sc_hd__a221o_1 _06910_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[13] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[13] ),
    .C1(net1243),
    .X(_02380_));
 sky130_fd_sc_hd__o22a_1 _06911_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[13] ),
    .A2(net1229),
    .B1(_02379_),
    .B2(_02380_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__nor2_1 _06912_ (.A(_00940_),
    .B(net1213),
    .Y(_02381_));
 sky130_fd_sc_hd__a221o_1 _06913_ (.A1(net1279),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[14] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[14] ),
    .C1(net1243),
    .X(_02382_));
 sky130_fd_sc_hd__o22a_1 _06914_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[14] ),
    .A2(net1229),
    .B1(_02381_),
    .B2(_02382_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__and3_1 _06915_ (.A(net1354),
    .B(net1261),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[15] ),
    .X(_02383_));
 sky130_fd_sc_hd__a221o_1 _06916_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[15] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ),
    .C1(net1245),
    .X(_02384_));
 sky130_fd_sc_hd__o22a_1 _06917_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[15] ),
    .A2(net1229),
    .B1(_02383_),
    .B2(_02384_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__and3_1 _06918_ (.A(net1360),
    .B(net1261),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[16] ),
    .X(_02385_));
 sky130_fd_sc_hd__a221o_1 _06919_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[16] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ),
    .C1(net1245),
    .X(_02386_));
 sky130_fd_sc_hd__o22a_1 _06920_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[16] ),
    .A2(net1233),
    .B1(_02385_),
    .B2(_02386_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__and3_1 _06921_ (.A(net1360),
    .B(net1368),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ),
    .X(_02387_));
 sky130_fd_sc_hd__a221o_1 _06922_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[17] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[17] ),
    .C1(net1245),
    .X(_02388_));
 sky130_fd_sc_hd__o22a_1 _06923_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[17] ),
    .A2(net1233),
    .B1(_02387_),
    .B2(_02388_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__and3_1 _06924_ (.A(net1360),
    .B(net1368),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ),
    .X(_02389_));
 sky130_fd_sc_hd__a221o_1 _06925_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[18] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[18] ),
    .C1(net1245),
    .X(_02390_));
 sky130_fd_sc_hd__o22a_1 _06926_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[18] ),
    .A2(net1230),
    .B1(_02389_),
    .B2(_02390_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__and3_1 _06927_ (.A(net1361),
    .B(net1265),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[19] ),
    .X(_02391_));
 sky130_fd_sc_hd__a221o_1 _06928_ (.A1(net1278),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[19] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ),
    .C1(net1245),
    .X(_02392_));
 sky130_fd_sc_hd__o22a_1 _06929_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[19] ),
    .A2(net1230),
    .B1(_02391_),
    .B2(_02392_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__and3_1 _06930_ (.A(net1359),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ),
    .X(_02393_));
 sky130_fd_sc_hd__a221o_1 _06931_ (.A1(net1276),
    .A2(net2295),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[20] ),
    .C1(net1245),
    .X(_02394_));
 sky130_fd_sc_hd__o22a_1 _06932_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[20] ),
    .A2(net1226),
    .B1(_02393_),
    .B2(_02394_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__and3_1 _06933_ (.A(net1359),
    .B(net1261),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[21] ),
    .X(_02395_));
 sky130_fd_sc_hd__a221o_1 _06934_ (.A1(net1276),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[21] ),
    .B1(net1147),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ),
    .C1(net1245),
    .X(_02396_));
 sky130_fd_sc_hd__o22a_1 _06935_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[21] ),
    .A2(net1226),
    .B1(_02395_),
    .B2(_02396_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__and3_1 _06936_ (.A(net1358),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ),
    .X(_02397_));
 sky130_fd_sc_hd__a221o_1 _06937_ (.A1(net1276),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[22] ),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[22] ),
    .C1(net1245),
    .X(_02398_));
 sky130_fd_sc_hd__o22a_1 _06938_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[22] ),
    .A2(net1226),
    .B1(_02397_),
    .B2(_02398_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__and3_1 _06939_ (.A(net1360),
    .B(net1368),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ),
    .X(_02399_));
 sky130_fd_sc_hd__a221o_1 _06940_ (.A1(net1276),
    .A2(net2340),
    .B1(net1162),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[23] ),
    .C1(net1245),
    .X(_02400_));
 sky130_fd_sc_hd__o22a_1 _06941_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[23] ),
    .A2(net1229),
    .B1(_02399_),
    .B2(_02400_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__and3_1 _06942_ (.A(net1358),
    .B(net1264),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[24] ),
    .X(_02401_));
 sky130_fd_sc_hd__a221o_1 _06943_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[24] ),
    .B1(net1151),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ),
    .C1(net1249),
    .X(_02402_));
 sky130_fd_sc_hd__o22a_1 _06944_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[24] ),
    .A2(net1226),
    .B1(_02401_),
    .B2(_02402_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__nor2_1 _06945_ (.A(_00941_),
    .B(net1213),
    .Y(_02403_));
 sky130_fd_sc_hd__a221o_1 _06946_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[25] ),
    .B1(net1165),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[25] ),
    .C1(net1248),
    .X(_02404_));
 sky130_fd_sc_hd__o22a_1 _06947_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[25] ),
    .A2(net1226),
    .B1(_02403_),
    .B2(_02404_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__and3_1 _06948_ (.A(net1358),
    .B(net1262),
    .C(\u_pwm.u_pwm_0.u_reg.reg_2[26] ),
    .X(_02405_));
 sky130_fd_sc_hd__a221o_1 _06949_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[26] ),
    .B1(net1145),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ),
    .C1(net1249),
    .X(_02406_));
 sky130_fd_sc_hd__o22a_1 _06950_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[26] ),
    .A2(net1226),
    .B1(_02405_),
    .B2(_02406_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__and3_1 _06951_ (.A(net1359),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .X(_02407_));
 sky130_fd_sc_hd__a221o_1 _06952_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[27] ),
    .B1(net1161),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[27] ),
    .C1(net1249),
    .X(_02408_));
 sky130_fd_sc_hd__o22a_1 _06953_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[27] ),
    .A2(net1226),
    .B1(_02407_),
    .B2(_02408_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__and3_1 _06954_ (.A(net1358),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ),
    .X(_02409_));
 sky130_fd_sc_hd__a221o_1 _06955_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[28] ),
    .B1(net1160),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[28] ),
    .C1(net1248),
    .X(_02410_));
 sky130_fd_sc_hd__o22a_1 _06956_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[28] ),
    .A2(net1227),
    .B1(_02409_),
    .B2(_02410_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__and3_1 _06957_ (.A(net1358),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ),
    .X(_02411_));
 sky130_fd_sc_hd__a221o_1 _06958_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[29] ),
    .B1(net1160),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[29] ),
    .C1(net1249),
    .X(_02412_));
 sky130_fd_sc_hd__o22a_1 _06959_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[29] ),
    .A2(net1227),
    .B1(_02411_),
    .B2(_02412_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__and3_1 _06960_ (.A(net1358),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .X(_02413_));
 sky130_fd_sc_hd__a221o_1 _06961_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[30] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[30] ),
    .C1(net1252),
    .X(_02414_));
 sky130_fd_sc_hd__o22a_1 _06962_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[30] ),
    .A2(net1227),
    .B1(_02413_),
    .B2(_02414_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__and3_1 _06963_ (.A(net1359),
    .B(net1365),
    .C(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ),
    .X(_02415_));
 sky130_fd_sc_hd__a221o_1 _06964_ (.A1(net1281),
    .A2(\u_pwm.u_pwm_0.u_reg.reg_1[31] ),
    .B1(net1163),
    .B2(\u_pwm.u_pwm_0.u_reg.reg_2[31] ),
    .C1(net1252),
    .X(_02416_));
 sky130_fd_sc_hd__o22a_1 _06965_ (.A1(\u_pwm.u_pwm_0.u_reg.reg_0[31] ),
    .A2(net1226),
    .B1(_02415_),
    .B2(_02416_),
    .X(\u_pwm.u_pwm_0.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__xnor2_4 _06966_ (.A(net1070),
    .B(net1073),
    .Y(_02417_));
 sky130_fd_sc_hd__xnor2_4 _06967_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .Y(_02418_));
 sky130_fd_sc_hd__o22a_1 _06968_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ),
    .A2(_02417_),
    .B1(_02418_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ),
    .X(_02419_));
 sky130_fd_sc_hd__xnor2_4 _06969_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .Y(_02420_));
 sky130_fd_sc_hd__xnor2_4 _06970_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ),
    .Y(_02421_));
 sky130_fd_sc_hd__xnor2_4 _06971_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .Y(_02422_));
 sky130_fd_sc_hd__xnor2_2 _06972_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ),
    .Y(_02423_));
 sky130_fd_sc_hd__o211a_1 _06973_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ),
    .A2(_02422_),
    .B1(_02423_),
    .C1(\u_pwm.u_pwm_2.cfg_pwm_comp2[0] ),
    .X(_02424_));
 sky130_fd_sc_hd__xnor2_4 _06974_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ),
    .Y(_02425_));
 sky130_fd_sc_hd__a221o_1 _06975_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ),
    .A2(_02422_),
    .B1(_02425_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ),
    .C1(_02424_),
    .X(_02426_));
 sky130_fd_sc_hd__xnor2_4 _06976_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ),
    .Y(_02427_));
 sky130_fd_sc_hd__o22a_1 _06977_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ),
    .A2(_02425_),
    .B1(_02427_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ),
    .X(_02428_));
 sky130_fd_sc_hd__xnor2_4 _06978_ (.A(net1071),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .Y(_02429_));
 sky130_fd_sc_hd__a22o_1 _06979_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ),
    .A2(_02427_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ),
    .X(_02430_));
 sky130_fd_sc_hd__a21o_1 _06980_ (.A1(_02426_),
    .A2(_02428_),
    .B1(_02430_),
    .X(_02431_));
 sky130_fd_sc_hd__o22a_1 _06981_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ),
    .A2(_02421_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ),
    .X(_02432_));
 sky130_fd_sc_hd__a22o_1 _06982_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ),
    .A2(_02420_),
    .B1(_02421_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ),
    .X(_02433_));
 sky130_fd_sc_hd__a21o_1 _06983_ (.A1(_02431_),
    .A2(_02432_),
    .B1(_02433_),
    .X(_02434_));
 sky130_fd_sc_hd__xnor2_4 _06984_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .Y(_02435_));
 sky130_fd_sc_hd__o22a_1 _06985_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ),
    .A2(_02420_),
    .B1(_02435_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ),
    .X(_02436_));
 sky130_fd_sc_hd__xnor2_4 _06986_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .Y(_02437_));
 sky130_fd_sc_hd__a22o_1 _06987_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ),
    .A2(_02435_),
    .B1(_02437_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ),
    .X(_02438_));
 sky130_fd_sc_hd__a21o_1 _06988_ (.A1(_02434_),
    .A2(_02436_),
    .B1(_02438_),
    .X(_02439_));
 sky130_fd_sc_hd__xnor2_4 _06989_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .Y(_02440_));
 sky130_fd_sc_hd__o221a_1 _06990_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ),
    .A2(_02437_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ),
    .C1(_02439_),
    .X(_02441_));
 sky130_fd_sc_hd__a221o_1 _06991_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ),
    .A2(_02417_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ),
    .C1(_02441_),
    .X(_02442_));
 sky130_fd_sc_hd__xnor2_4 _06992_ (.A(net1070),
    .B(net1072),
    .Y(_02443_));
 sky130_fd_sc_hd__o21bai_1 _06993_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .A2(_02443_),
    .B1_N(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ),
    .Y(_02444_));
 sky130_fd_sc_hd__a21o_1 _06994_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .A2(_02443_),
    .B1(_02444_),
    .X(_02445_));
 sky130_fd_sc_hd__xnor2_4 _06995_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .Y(_02446_));
 sky130_fd_sc_hd__xnor2_4 _06996_ (.A(net1070),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .Y(_02447_));
 sky130_fd_sc_hd__o22a_1 _06997_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ),
    .A2(_02446_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .X(_02448_));
 sky130_fd_sc_hd__inv_2 _06998_ (.A(_02448_),
    .Y(_02449_));
 sky130_fd_sc_hd__a211o_1 _06999_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ),
    .A2(_02446_),
    .B1(_02449_),
    .C1(_02445_),
    .X(_02450_));
 sky130_fd_sc_hd__a221o_1 _07000_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ),
    .A2(_02418_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .C1(_02450_),
    .X(_02451_));
 sky130_fd_sc_hd__a21o_1 _07001_ (.A1(_02419_),
    .A2(_02442_),
    .B1(_02451_),
    .X(_02452_));
 sky130_fd_sc_hd__a211o_1 _07002_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .A2(_02447_),
    .B1(_02448_),
    .C1(_02445_),
    .X(_02453_));
 sky130_fd_sc_hd__o311a_1 _07003_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .A3(_02443_),
    .B1(_02453_),
    .C1(\u_pwm.u_pwm_2.cfg_comp2_center ),
    .X(_02454_));
 sky130_fd_sc_hd__o211a_1 _07004_ (.A1(_00912_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[0] ),
    .C1(_00913_),
    .X(_02455_));
 sky130_fd_sc_hd__a221o_1 _07005_ (.A1(net725),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ),
    .B2(_00912_),
    .C1(_02455_),
    .X(_02456_));
 sky130_fd_sc_hd__o221a_1 _07006_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ),
    .B2(net725),
    .C1(_02456_),
    .X(_02457_));
 sky130_fd_sc_hd__a221o_1 _07007_ (.A1(_00909_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ),
    .B2(_00910_),
    .C1(_02457_),
    .X(_02458_));
 sky130_fd_sc_hd__o221a_1 _07008_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ),
    .B2(_00909_),
    .C1(_02458_),
    .X(_02459_));
 sky130_fd_sc_hd__a221o_1 _07009_ (.A1(_00907_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ),
    .B2(_00908_),
    .C1(_02459_),
    .X(_02460_));
 sky130_fd_sc_hd__o221a_1 _07010_ (.A1(_00906_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ),
    .B2(_00907_),
    .C1(_02460_),
    .X(_02461_));
 sky130_fd_sc_hd__o22a_1 _07011_ (.A1(_00900_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ),
    .B2(_00901_),
    .X(_02462_));
 sky130_fd_sc_hd__o22a_1 _07012_ (.A1(_00904_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ),
    .B2(_00905_),
    .X(_02463_));
 sky130_fd_sc_hd__o22a_1 _07013_ (.A1(_00902_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ),
    .B2(_00903_),
    .X(_02464_));
 sky130_fd_sc_hd__nand2_1 _07014_ (.A(_00900_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .Y(_02465_));
 sky130_fd_sc_hd__nand2_1 _07015_ (.A(_00899_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .Y(_02466_));
 sky130_fd_sc_hd__a22oi_1 _07016_ (.A1(_00901_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ),
    .B2(_00902_),
    .Y(_02467_));
 sky130_fd_sc_hd__a22oi_1 _07017_ (.A1(_00903_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ),
    .B2(_00904_),
    .Y(_02468_));
 sky130_fd_sc_hd__inv_2 _07018_ (.A(_02468_),
    .Y(_02469_));
 sky130_fd_sc_hd__nand2_1 _07019_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ),
    .Y(_02470_));
 sky130_fd_sc_hd__nor2_1 _07020_ (.A(_00899_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .Y(_02471_));
 sky130_fd_sc_hd__a221o_1 _07021_ (.A1(_00905_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ),
    .B2(_00906_),
    .C1(_02471_),
    .X(_02472_));
 sky130_fd_sc_hd__and2b_1 _07022_ (.A_N(_02472_),
    .B(_02470_),
    .X(_02473_));
 sky130_fd_sc_hd__and4_1 _07023_ (.A(_02463_),
    .B(_02464_),
    .C(_02467_),
    .D(_02468_),
    .X(_02474_));
 sky130_fd_sc_hd__and3_1 _07024_ (.A(_02462_),
    .B(_02465_),
    .C(_02466_),
    .X(_02475_));
 sky130_fd_sc_hd__and4b_1 _07025_ (.A_N(_02461_),
    .B(_02473_),
    .C(_02474_),
    .D(_02475_),
    .X(_02476_));
 sky130_fd_sc_hd__o21ai_1 _07026_ (.A1(_02463_),
    .A2(_02469_),
    .B1(_02464_),
    .Y(_02477_));
 sky130_fd_sc_hd__a21bo_1 _07027_ (.A1(_02467_),
    .A2(_02477_),
    .B1_N(_02462_),
    .X(_02478_));
 sky130_fd_sc_hd__a31o_1 _07028_ (.A1(_02465_),
    .A2(_02466_),
    .A3(_02478_),
    .B1(_02471_),
    .X(_02479_));
 sky130_fd_sc_hd__nor2_1 _07029_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ),
    .Y(_02480_));
 sky130_fd_sc_hd__a211o_1 _07030_ (.A1(_02470_),
    .A2(_02479_),
    .B1(_02480_),
    .C1(\u_pwm.u_pwm_2.cfg_comp2_center ),
    .X(_02481_));
 sky130_fd_sc_hd__o2bb2a_1 _07031_ (.A1_N(_02452_),
    .A2_N(_02454_),
    .B1(_02476_),
    .B2(_02481_),
    .X(_02482_));
 sky130_fd_sc_hd__o22a_1 _07032_ (.A1(_00904_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[9] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[8] ),
    .B2(_00905_),
    .X(_02483_));
 sky130_fd_sc_hd__nand2b_1 _07033_ (.A_N(\u_pwm.u_pwm_2.cfg_pwm_comp0[1] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .Y(_02484_));
 sky130_fd_sc_hd__and2b_1 _07034_ (.A_N(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp0[2] ),
    .X(_02485_));
 sky130_fd_sc_hd__and2b_1 _07035_ (.A_N(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp0[1] ),
    .X(_02486_));
 sky130_fd_sc_hd__a311o_1 _07036_ (.A1(_00913_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[0] ),
    .A3(_02484_),
    .B1(_02485_),
    .C1(_02486_),
    .X(_02487_));
 sky130_fd_sc_hd__o22a_1 _07037_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[3] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[2] ),
    .B2(net725),
    .X(_02488_));
 sky130_fd_sc_hd__a22o_1 _07038_ (.A1(_00909_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[4] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[3] ),
    .B2(_00910_),
    .X(_02489_));
 sky130_fd_sc_hd__a21o_1 _07039_ (.A1(_02487_),
    .A2(_02488_),
    .B1(_02489_),
    .X(_02490_));
 sky130_fd_sc_hd__o22a_1 _07040_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[4] ),
    .B2(_00909_),
    .X(_02491_));
 sky130_fd_sc_hd__a22o_1 _07041_ (.A1(_00907_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ),
    .B2(_00908_),
    .X(_02492_));
 sky130_fd_sc_hd__a21o_1 _07042_ (.A1(_02490_),
    .A2(_02491_),
    .B1(_02492_),
    .X(_02493_));
 sky130_fd_sc_hd__o221a_1 _07043_ (.A1(_00906_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ),
    .B2(_00907_),
    .C1(_02493_),
    .X(_02494_));
 sky130_fd_sc_hd__a22o_1 _07044_ (.A1(_00905_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[8] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ),
    .B2(_00906_),
    .X(_02495_));
 sky130_fd_sc_hd__o21ai_1 _07045_ (.A1(_02494_),
    .A2(_02495_),
    .B1(_02483_),
    .Y(_02496_));
 sky130_fd_sc_hd__o2bb2a_1 _07046_ (.A1_N(\u_pwm.u_pwm_2.cfg_pwm_comp0[9] ),
    .A2_N(_00904_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[10] ),
    .B2(_00945_),
    .X(_02497_));
 sky130_fd_sc_hd__a2bb2o_1 _07047_ (.A1_N(_00902_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ),
    .B1(_00945_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[10] ),
    .X(_02498_));
 sky130_fd_sc_hd__a21oi_1 _07048_ (.A1(_02496_),
    .A2(_02497_),
    .B1(_02498_),
    .Y(_02499_));
 sky130_fd_sc_hd__a2bb2o_1 _07049_ (.A1_N(_00898_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_comp0[15] ),
    .B1(_00943_),
    .B2(net1072),
    .X(_02500_));
 sky130_fd_sc_hd__nand2_1 _07050_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp0[15] ),
    .Y(_02501_));
 sky130_fd_sc_hd__nor2_1 _07051_ (.A(net1072),
    .B(_00943_),
    .Y(_02502_));
 sky130_fd_sc_hd__or3b_1 _07052_ (.A(_02502_),
    .B(_02500_),
    .C_N(_02501_),
    .X(_02503_));
 sky130_fd_sc_hd__a2bb2o_1 _07053_ (.A1_N(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ),
    .A2_N(_00901_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .B2(_00944_),
    .X(_02504_));
 sky130_fd_sc_hd__nor2_1 _07054_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .B(_00944_),
    .Y(_02505_));
 sky130_fd_sc_hd__a221o_1 _07055_ (.A1(_00901_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ),
    .B2(_00902_),
    .C1(_02505_),
    .X(_02506_));
 sky130_fd_sc_hd__or4_1 _07056_ (.A(_02499_),
    .B(_02503_),
    .C(_02504_),
    .D(_02506_),
    .X(_02507_));
 sky130_fd_sc_hd__or3b_1 _07057_ (.A(_02505_),
    .B(_02503_),
    .C_N(_02504_),
    .X(_02508_));
 sky130_fd_sc_hd__a21oi_1 _07058_ (.A1(_02500_),
    .A2(_02501_),
    .B1(\u_pwm.u_pwm_2.cfg_comp0_center ),
    .Y(_02509_));
 sky130_fd_sc_hd__o22a_1 _07059_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[14] ),
    .A2(_02443_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[13] ),
    .X(_02510_));
 sky130_fd_sc_hd__nor2_1 _07060_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ),
    .B(_02446_),
    .Y(_02511_));
 sky130_fd_sc_hd__o22a_1 _07061_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[10] ),
    .A2(_02417_),
    .B1(_02418_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ),
    .X(_02512_));
 sky130_fd_sc_hd__a22o_1 _07062_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[10] ),
    .A2(_02417_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[9] ),
    .X(_02513_));
 sky130_fd_sc_hd__o22a_1 _07063_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[8] ),
    .A2(_02437_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[9] ),
    .X(_02514_));
 sky130_fd_sc_hd__or2_1 _07064_ (.A(_02513_),
    .B(_02514_),
    .X(_02515_));
 sky130_fd_sc_hd__a22o_1 _07065_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ),
    .A2(_02418_),
    .B1(_02512_),
    .B2(_02515_),
    .X(_02516_));
 sky130_fd_sc_hd__o211a_1 _07066_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[1] ),
    .A2(_02422_),
    .B1(_02423_),
    .C1(\u_pwm.u_pwm_2.cfg_pwm_comp0[0] ),
    .X(_02517_));
 sky130_fd_sc_hd__a22o_1 _07067_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[1] ),
    .A2(_02422_),
    .B1(_02425_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[2] ),
    .X(_02518_));
 sky130_fd_sc_hd__o22a_1 _07068_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[2] ),
    .A2(_02425_),
    .B1(_02427_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[3] ),
    .X(_02519_));
 sky130_fd_sc_hd__o21a_1 _07069_ (.A1(_02517_),
    .A2(_02518_),
    .B1(_02519_),
    .X(_02520_));
 sky130_fd_sc_hd__a22o_1 _07070_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[3] ),
    .A2(_02427_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[4] ),
    .X(_02521_));
 sky130_fd_sc_hd__o22a_1 _07071_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ),
    .A2(_02421_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[4] ),
    .X(_02522_));
 sky130_fd_sc_hd__o21a_1 _07072_ (.A1(_02520_),
    .A2(_02521_),
    .B1(_02522_),
    .X(_02523_));
 sky130_fd_sc_hd__a22o_1 _07073_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ),
    .A2(_02420_),
    .B1(_02421_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ),
    .X(_02524_));
 sky130_fd_sc_hd__or2_1 _07074_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ),
    .B(_02435_),
    .X(_02525_));
 sky130_fd_sc_hd__o221a_1 _07075_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ),
    .A2(_02420_),
    .B1(_02523_),
    .B2(_02524_),
    .C1(_02525_),
    .X(_02526_));
 sky130_fd_sc_hd__a22o_1 _07076_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ),
    .A2(_02418_),
    .B1(_02437_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[8] ),
    .X(_02527_));
 sky130_fd_sc_hd__a211o_1 _07077_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ),
    .A2(_02435_),
    .B1(_02511_),
    .C1(_02527_),
    .X(_02528_));
 sky130_fd_sc_hd__nand2_1 _07078_ (.A(_02512_),
    .B(_02514_),
    .Y(_02529_));
 sky130_fd_sc_hd__or3_1 _07079_ (.A(_02513_),
    .B(_02528_),
    .C(_02529_),
    .X(_02530_));
 sky130_fd_sc_hd__o221a_1 _07080_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ),
    .A2(_02446_),
    .B1(_02526_),
    .B2(_02530_),
    .C1(_02516_),
    .X(_02531_));
 sky130_fd_sc_hd__a221o_1 _07081_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ),
    .A2(_02446_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp0[13] ),
    .C1(_02531_),
    .X(_02532_));
 sky130_fd_sc_hd__a221o_1 _07082_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp0[14] ),
    .A2(_02443_),
    .B1(_02510_),
    .B2(_02532_),
    .C1(\u_pwm.u_pwm_2.cfg_pwm_comp0[15] ),
    .X(_02533_));
 sky130_fd_sc_hd__a32o_1 _07083_ (.A1(_02507_),
    .A2(_02508_),
    .A3(_02509_),
    .B1(_02533_),
    .B2(\u_pwm.u_pwm_2.cfg_comp0_center ),
    .X(_02534_));
 sky130_fd_sc_hd__inv_2 _07084_ (.A(_02534_),
    .Y(_02535_));
 sky130_fd_sc_hd__o22a_1 _07085_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[12] ),
    .A2(_02446_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[13] ),
    .X(_02536_));
 sky130_fd_sc_hd__a22oi_1 _07086_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[11] ),
    .A2(_02418_),
    .B1(_02446_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[12] ),
    .Y(_02537_));
 sky130_fd_sc_hd__o22a_1 _07087_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[10] ),
    .A2(_02417_),
    .B1(_02418_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[11] ),
    .X(_02538_));
 sky130_fd_sc_hd__a22o_1 _07088_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[10] ),
    .A2(_02417_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[9] ),
    .X(_02539_));
 sky130_fd_sc_hd__o22a_1 _07089_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[8] ),
    .A2(_02437_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[9] ),
    .X(_02540_));
 sky130_fd_sc_hd__o211a_1 _07090_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[1] ),
    .A2(_02422_),
    .B1(_02423_),
    .C1(\u_pwm.u_pwm_2.cfg_pwm_comp1[0] ),
    .X(_02541_));
 sky130_fd_sc_hd__a22o_1 _07091_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[1] ),
    .A2(_02422_),
    .B1(_02425_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[2] ),
    .X(_02542_));
 sky130_fd_sc_hd__or2_1 _07092_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[2] ),
    .B(_02425_),
    .X(_02543_));
 sky130_fd_sc_hd__o221a_1 _07093_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[3] ),
    .A2(_02427_),
    .B1(_02541_),
    .B2(_02542_),
    .C1(_02543_),
    .X(_02544_));
 sky130_fd_sc_hd__a22o_1 _07094_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[3] ),
    .A2(_02427_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[4] ),
    .X(_02545_));
 sky130_fd_sc_hd__o22a_1 _07095_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[5] ),
    .A2(_02421_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[4] ),
    .X(_02546_));
 sky130_fd_sc_hd__o21a_1 _07096_ (.A1(_02544_),
    .A2(_02545_),
    .B1(_02546_),
    .X(_02547_));
 sky130_fd_sc_hd__a221o_1 _07097_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[6] ),
    .A2(_02420_),
    .B1(_02421_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[5] ),
    .C1(_02547_),
    .X(_02548_));
 sky130_fd_sc_hd__o22a_1 _07098_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[6] ),
    .A2(_02420_),
    .B1(_02435_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[7] ),
    .X(_02549_));
 sky130_fd_sc_hd__o21ai_1 _07099_ (.A1(_02539_),
    .A2(_02540_),
    .B1(_02538_),
    .Y(_02550_));
 sky130_fd_sc_hd__nand2_1 _07100_ (.A(_02537_),
    .B(_02550_),
    .Y(_02551_));
 sky130_fd_sc_hd__a221o_1 _07101_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[7] ),
    .A2(_02435_),
    .B1(_02437_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[8] ),
    .C1(_02539_),
    .X(_02552_));
 sky130_fd_sc_hd__nand4_1 _07102_ (.A(_02536_),
    .B(_02537_),
    .C(_02538_),
    .D(_02540_),
    .Y(_02553_));
 sky130_fd_sc_hd__a211o_1 _07103_ (.A1(_02548_),
    .A2(_02549_),
    .B1(_02552_),
    .C1(_02553_),
    .X(_02554_));
 sky130_fd_sc_hd__xnor2_1 _07104_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[14] ),
    .B(_02443_),
    .Y(_02555_));
 sky130_fd_sc_hd__a32o_1 _07105_ (.A1(_02536_),
    .A2(_02551_),
    .A3(_02554_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp1[13] ),
    .X(_02556_));
 sky130_fd_sc_hd__or3_1 _07106_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp1[15] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp1[14] ),
    .C(_02443_),
    .X(_02557_));
 sky130_fd_sc_hd__o311a_1 _07107_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp1[15] ),
    .A2(_02555_),
    .A3(_02556_),
    .B1(_02557_),
    .C1(\u_pwm.u_pwm_2.cfg_comp1_center ),
    .X(_02558_));
 sky130_fd_sc_hd__a2bb2o_1 _07108_ (.A1_N(_00902_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_comp1[11] ),
    .B1(_00947_),
    .B2(net1073),
    .X(_02559_));
 sky130_fd_sc_hd__a22o_1 _07109_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .A2(_00950_),
    .B1(_00951_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .X(_02560_));
 sky130_fd_sc_hd__o211a_1 _07110_ (.A1(_00912_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[1] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[0] ),
    .C1(_00913_),
    .X(_02561_));
 sky130_fd_sc_hd__a22o_1 _07111_ (.A1(net725),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[2] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[1] ),
    .B2(_00912_),
    .X(_02562_));
 sky130_fd_sc_hd__o22a_1 _07112_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[3] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[2] ),
    .B2(net725),
    .X(_02563_));
 sky130_fd_sc_hd__o21ai_1 _07113_ (.A1(_02561_),
    .A2(_02562_),
    .B1(_02563_),
    .Y(_02564_));
 sky130_fd_sc_hd__a22oi_1 _07114_ (.A1(_00909_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[4] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[3] ),
    .B2(_00910_),
    .Y(_02565_));
 sky130_fd_sc_hd__o22a_1 _07115_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[5] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[4] ),
    .B2(_00909_),
    .X(_02566_));
 sky130_fd_sc_hd__a21bo_1 _07116_ (.A1(_02564_),
    .A2(_02565_),
    .B1_N(_02566_),
    .X(_02567_));
 sky130_fd_sc_hd__o2bb2a_1 _07117_ (.A1_N(\u_pwm.u_pwm_2.cfg_pwm_comp1[5] ),
    .A2_N(_00908_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .B2(_00951_),
    .X(_02568_));
 sky130_fd_sc_hd__a21o_1 _07118_ (.A1(_02567_),
    .A2(_02568_),
    .B1(_02560_),
    .X(_02569_));
 sky130_fd_sc_hd__o22a_1 _07119_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .A2(_00949_),
    .B1(_00950_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .X(_02570_));
 sky130_fd_sc_hd__a22o_1 _07120_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .A2(_00948_),
    .B1(_00949_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .X(_02571_));
 sky130_fd_sc_hd__a21o_1 _07121_ (.A1(_02569_),
    .A2(_02570_),
    .B1(_02571_),
    .X(_02572_));
 sky130_fd_sc_hd__o221a_1 _07122_ (.A1(net1073),
    .A2(_00947_),
    .B1(_00948_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .C1(_02572_),
    .X(_02573_));
 sky130_fd_sc_hd__o22a_1 _07123_ (.A1(_00898_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[15] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[14] ),
    .B2(_00899_),
    .X(_02574_));
 sky130_fd_sc_hd__nand2_1 _07124_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp1[15] ),
    .Y(_02575_));
 sky130_fd_sc_hd__o211a_1 _07125_ (.A1(net1072),
    .A2(_00946_),
    .B1(_02574_),
    .C1(_02575_),
    .X(_02576_));
 sky130_fd_sc_hd__o22ai_1 _07126_ (.A1(_00900_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp1[13] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp1[12] ),
    .B2(_00901_),
    .Y(_02577_));
 sky130_fd_sc_hd__nand2_1 _07127_ (.A(_00901_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp1[12] ),
    .Y(_02578_));
 sky130_fd_sc_hd__nand2_1 _07128_ (.A(_00900_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp1[13] ),
    .Y(_02579_));
 sky130_fd_sc_hd__nand2_1 _07129_ (.A(_00902_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp1[11] ),
    .Y(_02580_));
 sky130_fd_sc_hd__and3b_1 _07130_ (.A_N(_02577_),
    .B(_02578_),
    .C(_02579_),
    .X(_02581_));
 sky130_fd_sc_hd__o2111a_1 _07131_ (.A1(_02559_),
    .A2(_02573_),
    .B1(_02576_),
    .C1(_02580_),
    .D1(_02581_),
    .X(_02582_));
 sky130_fd_sc_hd__and2b_1 _07132_ (.A_N(_02574_),
    .B(_02575_),
    .X(_02583_));
 sky130_fd_sc_hd__a311o_1 _07133_ (.A1(_02576_),
    .A2(_02577_),
    .A3(_02579_),
    .B1(_02583_),
    .C1(\u_pwm.u_pwm_2.cfg_comp1_center ),
    .X(_02584_));
 sky130_fd_sc_hd__o21ba_1 _07134_ (.A1(_02582_),
    .A2(_02584_),
    .B1_N(_02558_),
    .X(_02585_));
 sky130_fd_sc_hd__xnor2_1 _07135_ (.A(_02534_),
    .B(_02585_),
    .Y(_02586_));
 sky130_fd_sc_hd__xnor2_1 _07136_ (.A(_02482_),
    .B(_02586_),
    .Y(_02587_));
 sky130_fd_sc_hd__o22a_1 _07137_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[10] ),
    .A2(_02417_),
    .B1(_02418_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .X(_02588_));
 sky130_fd_sc_hd__a22o_1 _07138_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[10] ),
    .A2(_02417_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[9] ),
    .X(_02589_));
 sky130_fd_sc_hd__o22a_1 _07139_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ),
    .A2(_02437_),
    .B1(_02440_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[9] ),
    .X(_02590_));
 sky130_fd_sc_hd__or2_1 _07140_ (.A(_02589_),
    .B(_02590_),
    .X(_02591_));
 sky130_fd_sc_hd__a22o_1 _07141_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .A2(_02418_),
    .B1(_02588_),
    .B2(_02591_),
    .X(_02592_));
 sky130_fd_sc_hd__o211a_1 _07142_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ),
    .A2(_02422_),
    .B1(_02423_),
    .C1(\u_pwm.u_pwm_2.cfg_pwm_comp3[0] ),
    .X(_02593_));
 sky130_fd_sc_hd__a22o_1 _07143_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ),
    .A2(_02422_),
    .B1(_02425_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ),
    .X(_02594_));
 sky130_fd_sc_hd__o22a_1 _07144_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ),
    .A2(_02425_),
    .B1(_02427_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ),
    .X(_02595_));
 sky130_fd_sc_hd__o21a_1 _07145_ (.A1(_02593_),
    .A2(_02594_),
    .B1(_02595_),
    .X(_02596_));
 sky130_fd_sc_hd__a22o_1 _07146_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ),
    .A2(_02427_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ),
    .X(_02597_));
 sky130_fd_sc_hd__o22a_1 _07147_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ),
    .A2(_02421_),
    .B1(_02429_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ),
    .X(_02598_));
 sky130_fd_sc_hd__o21a_1 _07148_ (.A1(_02596_),
    .A2(_02597_),
    .B1(_02598_),
    .X(_02599_));
 sky130_fd_sc_hd__a221o_1 _07149_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ),
    .A2(_02420_),
    .B1(_02421_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ),
    .C1(_02599_),
    .X(_02600_));
 sky130_fd_sc_hd__o221a_1 _07150_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ),
    .A2(_02420_),
    .B1(_02435_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ),
    .C1(_02600_),
    .X(_02601_));
 sky130_fd_sc_hd__a22o_1 _07151_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .A2(_02418_),
    .B1(_02435_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ),
    .X(_02602_));
 sky130_fd_sc_hd__a211o_1 _07152_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ),
    .A2(_02437_),
    .B1(_02589_),
    .C1(_02602_),
    .X(_02603_));
 sky130_fd_sc_hd__or4bb_1 _07153_ (.A(_02601_),
    .B(_02603_),
    .C_N(_02588_),
    .D_N(_02590_),
    .X(_02604_));
 sky130_fd_sc_hd__a22o_1 _07154_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ),
    .A2(_02446_),
    .B1(_02592_),
    .B2(_02604_),
    .X(_02605_));
 sky130_fd_sc_hd__o221a_1 _07155_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ),
    .A2(_02446_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[13] ),
    .C1(_02605_),
    .X(_02606_));
 sky130_fd_sc_hd__nor2_1 _07156_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ),
    .B(_02443_),
    .Y(_02607_));
 sky130_fd_sc_hd__a22o_1 _07157_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ),
    .A2(_02443_),
    .B1(_02447_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[13] ),
    .X(_02608_));
 sky130_fd_sc_hd__or4_1 _07158_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ),
    .B(_02606_),
    .C(_02607_),
    .D(_02608_),
    .X(_02609_));
 sky130_fd_sc_hd__or3_1 _07159_ (.A(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ),
    .C(_02443_),
    .X(_02610_));
 sky130_fd_sc_hd__and2_1 _07160_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ),
    .X(_02611_));
 sky130_fd_sc_hd__o22a_1 _07161_ (.A1(net1072),
    .A2(_00955_),
    .B1(_00956_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .X(_02612_));
 sky130_fd_sc_hd__a2bb2o_1 _07162_ (.A1_N(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ),
    .A2_N(_00901_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .B2(_00956_),
    .X(_02613_));
 sky130_fd_sc_hd__o22a_1 _07163_ (.A1(net1073),
    .A2(_00957_),
    .B1(_00958_),
    .B2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .X(_02614_));
 sky130_fd_sc_hd__a2bb2o_1 _07164_ (.A1_N(_00902_),
    .A2_N(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .B1(_00957_),
    .B2(net1073),
    .X(_02615_));
 sky130_fd_sc_hd__nand2_1 _07165_ (.A(_00901_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ),
    .Y(_02616_));
 sky130_fd_sc_hd__nand2_1 _07166_ (.A(_00902_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .Y(_02617_));
 sky130_fd_sc_hd__nand2_1 _07167_ (.A(_02616_),
    .B(_02617_),
    .Y(_02618_));
 sky130_fd_sc_hd__a2bb2o_1 _07168_ (.A1_N(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ),
    .A2_N(_00905_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .B2(_00958_),
    .X(_02619_));
 sky130_fd_sc_hd__a21o_1 _07169_ (.A1(_02614_),
    .A2(_02619_),
    .B1(_02615_),
    .X(_02620_));
 sky130_fd_sc_hd__a31o_1 _07170_ (.A1(_02616_),
    .A2(_02617_),
    .A3(_02620_),
    .B1(_02613_),
    .X(_02621_));
 sky130_fd_sc_hd__o2bb2a_1 _07171_ (.A1_N(_02621_),
    .A2_N(_02612_),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ),
    .B2(_00899_),
    .X(_02622_));
 sky130_fd_sc_hd__o211a_1 _07172_ (.A1(_00912_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[0] ),
    .C1(_00913_),
    .X(_02623_));
 sky130_fd_sc_hd__a221o_1 _07173_ (.A1(net725),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ),
    .B2(_00912_),
    .C1(_02623_),
    .X(_02624_));
 sky130_fd_sc_hd__o221a_1 _07174_ (.A1(_00910_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ),
    .B2(net725),
    .C1(_02624_),
    .X(_02625_));
 sky130_fd_sc_hd__a221o_1 _07175_ (.A1(_00909_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ),
    .B2(_00910_),
    .C1(_02625_),
    .X(_02626_));
 sky130_fd_sc_hd__o221a_1 _07176_ (.A1(_00908_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ),
    .B2(_00909_),
    .C1(_02626_),
    .X(_02627_));
 sky130_fd_sc_hd__a221o_1 _07177_ (.A1(_00907_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ),
    .B2(_00908_),
    .C1(_02627_),
    .X(_02628_));
 sky130_fd_sc_hd__o221a_1 _07178_ (.A1(_00906_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ),
    .B2(_00907_),
    .C1(_02628_),
    .X(_02629_));
 sky130_fd_sc_hd__nand2b_1 _07179_ (.A_N(_02613_),
    .B(_02614_),
    .Y(_02630_));
 sky130_fd_sc_hd__a221o_1 _07180_ (.A1(_00905_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ),
    .B1(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ),
    .B2(_00906_),
    .C1(_02611_),
    .X(_02631_));
 sky130_fd_sc_hd__nor2_1 _07181_ (.A(_00898_),
    .B(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ),
    .Y(_02632_));
 sky130_fd_sc_hd__a211o_1 _07182_ (.A1(net1072),
    .A2(_00955_),
    .B1(_02618_),
    .C1(_02632_),
    .X(_02633_));
 sky130_fd_sc_hd__or4_1 _07183_ (.A(_02615_),
    .B(_02619_),
    .C(_02631_),
    .D(_02633_),
    .X(_02634_));
 sky130_fd_sc_hd__or4b_1 _07184_ (.A(_02629_),
    .B(_02630_),
    .C(_02634_),
    .D_N(_02612_),
    .X(_02635_));
 sky130_fd_sc_hd__nor2_1 _07185_ (.A(\u_pwm.u_pwm_2.cfg_comp3_center ),
    .B(_02632_),
    .Y(_02636_));
 sky130_fd_sc_hd__o211a_1 _07186_ (.A1(_02611_),
    .A2(_02622_),
    .B1(_02635_),
    .C1(_02636_),
    .X(_02637_));
 sky130_fd_sc_hd__a31o_1 _07187_ (.A1(\u_pwm.u_pwm_2.cfg_comp3_center ),
    .A2(_02609_),
    .A3(_02610_),
    .B1(_02637_),
    .X(_02638_));
 sky130_fd_sc_hd__nand2_1 _07188_ (.A(_02587_),
    .B(_02638_),
    .Y(_02639_));
 sky130_fd_sc_hd__or2_1 _07189_ (.A(_02587_),
    .B(_02638_),
    .X(_02640_));
 sky130_fd_sc_hd__and4_1 _07190_ (.A(\u_pwm.u_pwm_2.cfg_pwm_mode[1] ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_mode[0] ),
    .C(_02639_),
    .D(_02640_),
    .X(_02641_));
 sky130_fd_sc_hd__nand2b_1 _07191_ (.A_N(\u_pwm.u_pwm_2.cfg_pwm_mode[1] ),
    .B(_02586_),
    .Y(_02642_));
 sky130_fd_sc_hd__a22oi_1 _07192_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_mode[1] ),
    .A2(_02587_),
    .B1(_02642_),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_mode[0] ),
    .Y(_02643_));
 sky130_fd_sc_hd__o32a_1 _07193_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_mode[1] ),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_mode[0] ),
    .A3(_02535_),
    .B1(_02641_),
    .B2(_02643_),
    .X(\u_pwm.u_pwm_2.u_pwm.pwm_wfm_i ));
 sky130_fd_sc_hd__and3_1 _07194_ (.A(net1350),
    .B(net1363),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[0] ),
    .X(_02644_));
 sky130_fd_sc_hd__a221o_1 _07195_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[0] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[0] ),
    .C1(net1236),
    .X(_02645_));
 sky130_fd_sc_hd__o22a_1 _07196_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[0] ),
    .A2(net1220),
    .B1(_02644_),
    .B2(_02645_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__and3_1 _07197_ (.A(net1350),
    .B(net1363),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ),
    .X(_02646_));
 sky130_fd_sc_hd__a221o_1 _07198_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[1] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[1] ),
    .C1(net1238),
    .X(_02647_));
 sky130_fd_sc_hd__o22a_1 _07199_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[1] ),
    .A2(net1220),
    .B1(_02646_),
    .B2(_02647_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__nor2_1 _07200_ (.A(_00954_),
    .B(net1211),
    .Y(_02648_));
 sky130_fd_sc_hd__a221o_1 _07201_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[2] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[2] ),
    .C1(net1238),
    .X(_02649_));
 sky130_fd_sc_hd__o22a_1 _07202_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[2] ),
    .A2(net1220),
    .B1(_02648_),
    .B2(_02649_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__and3_1 _07203_ (.A(net1351),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[3] ),
    .X(_02650_));
 sky130_fd_sc_hd__a221o_1 _07204_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[3] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ),
    .C1(net1238),
    .X(_02651_));
 sky130_fd_sc_hd__o22a_1 _07205_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[3] ),
    .A2(net1220),
    .B1(_02650_),
    .B2(_02651_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__and3_1 _07206_ (.A(net1350),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[4] ),
    .X(_02652_));
 sky130_fd_sc_hd__a221o_1 _07207_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[4] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ),
    .C1(net1236),
    .X(_02653_));
 sky130_fd_sc_hd__o22a_1 _07208_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[4] ),
    .A2(net1219),
    .B1(_02652_),
    .B2(_02653_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__nor2_1 _07209_ (.A(_00953_),
    .B(net1211),
    .Y(_02654_));
 sky130_fd_sc_hd__a221o_1 _07210_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[5] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[5] ),
    .C1(net1236),
    .X(_02655_));
 sky130_fd_sc_hd__o22a_1 _07211_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[5] ),
    .A2(net1219),
    .B1(_02654_),
    .B2(_02655_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__and3_1 _07212_ (.A(net1350),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[6] ),
    .X(_02656_));
 sky130_fd_sc_hd__a221o_1 _07213_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[6] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ),
    .C1(net1236),
    .X(_02657_));
 sky130_fd_sc_hd__o22a_1 _07214_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[6] ),
    .A2(net1219),
    .B1(_02656_),
    .B2(_02657_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__nor2_1 _07215_ (.A(_00952_),
    .B(net1211),
    .Y(_02658_));
 sky130_fd_sc_hd__a221o_1 _07216_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[7] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[7] ),
    .C1(net1238),
    .X(_02659_));
 sky130_fd_sc_hd__o22a_1 _07217_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[7] ),
    .A2(net1219),
    .B1(_02658_),
    .B2(_02659_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__and3_1 _07218_ (.A(net1349),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ),
    .X(_02660_));
 sky130_fd_sc_hd__a221o_1 _07219_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[8] ),
    .B1(net1156),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[8] ),
    .C1(net1237),
    .X(_02661_));
 sky130_fd_sc_hd__o22a_1 _07220_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[8] ),
    .A2(net1218),
    .B1(_02660_),
    .B2(_02661_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__and3_1 _07221_ (.A(net1349),
    .B(net1257),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[9] ),
    .X(_02662_));
 sky130_fd_sc_hd__a221o_1 _07222_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[9] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ),
    .C1(net1235),
    .X(_02663_));
 sky130_fd_sc_hd__o22a_1 _07223_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[9] ),
    .A2(net1218),
    .B1(_02662_),
    .B2(_02663_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__and3_1 _07224_ (.A(net1349),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ),
    .X(_02664_));
 sky130_fd_sc_hd__a221o_1 _07225_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[10] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[10] ),
    .C1(net1235),
    .X(_02665_));
 sky130_fd_sc_hd__o22a_1 _07226_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[10] ),
    .A2(net1218),
    .B1(_02664_),
    .B2(_02665_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__and3_1 _07227_ (.A(net1349),
    .B(net1257),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[11] ),
    .X(_02666_));
 sky130_fd_sc_hd__a221o_1 _07228_ (.A1(net1270),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[11] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ),
    .C1(net1235),
    .X(_02667_));
 sky130_fd_sc_hd__o22a_1 _07229_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[11] ),
    .A2(net1218),
    .B1(_02666_),
    .B2(_02667_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__and3_1 _07230_ (.A(net1348),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ),
    .X(_02668_));
 sky130_fd_sc_hd__a221o_1 _07231_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[12] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[12] ),
    .C1(net1234),
    .X(_02669_));
 sky130_fd_sc_hd__o22a_1 _07232_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[12] ),
    .A2(net1217),
    .B1(_02668_),
    .B2(_02669_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__and3_1 _07233_ (.A(net1348),
    .B(net1257),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[13] ),
    .X(_02670_));
 sky130_fd_sc_hd__a221o_1 _07234_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[13] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ),
    .C1(net1234),
    .X(_02671_));
 sky130_fd_sc_hd__o22a_1 _07235_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[13] ),
    .A2(net1218),
    .B1(_02670_),
    .B2(_02671_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__and3_1 _07236_ (.A(net1349),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ),
    .X(_02672_));
 sky130_fd_sc_hd__a221o_1 _07237_ (.A1(net1270),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[14] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[14] ),
    .C1(net1235),
    .X(_02673_));
 sky130_fd_sc_hd__o22a_1 _07238_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[14] ),
    .A2(net1218),
    .B1(_02672_),
    .B2(_02673_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__and3_1 _07239_ (.A(net1348),
    .B(net1257),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[15] ),
    .X(_02674_));
 sky130_fd_sc_hd__a221o_1 _07240_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[15] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ),
    .C1(net1235),
    .X(_02675_));
 sky130_fd_sc_hd__o22a_1 _07241_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[15] ),
    .A2(net1218),
    .B1(_02674_),
    .B2(_02675_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__and3_1 _07242_ (.A(net1350),
    .B(net1363),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[0] ),
    .X(_02676_));
 sky130_fd_sc_hd__a221o_1 _07243_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[16] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[16] ),
    .C1(net1236),
    .X(_02677_));
 sky130_fd_sc_hd__o22a_1 _07244_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[16] ),
    .A2(net1219),
    .B1(_02676_),
    .B2(_02677_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__and3_1 _07245_ (.A(net1350),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[17] ),
    .X(_02678_));
 sky130_fd_sc_hd__a221o_1 _07246_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[17] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ),
    .C1(net1236),
    .X(_02679_));
 sky130_fd_sc_hd__o22a_1 _07247_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[17] ),
    .A2(net1219),
    .B1(_02678_),
    .B2(_02679_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__and3_1 _07248_ (.A(net1350),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[18] ),
    .X(_02680_));
 sky130_fd_sc_hd__a221o_1 _07249_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[18] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ),
    .C1(net1236),
    .X(_02681_));
 sky130_fd_sc_hd__o22a_1 _07250_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[18] ),
    .A2(net1219),
    .B1(_02680_),
    .B2(_02681_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__and3_1 _07251_ (.A(net1350),
    .B(net1363),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ),
    .X(_02682_));
 sky130_fd_sc_hd__a221o_1 _07252_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[19] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[19] ),
    .C1(net1236),
    .X(_02683_));
 sky130_fd_sc_hd__o22a_1 _07253_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[19] ),
    .A2(net1219),
    .B1(_02682_),
    .B2(_02683_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__and3_1 _07254_ (.A(net1350),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[20] ),
    .X(_02684_));
 sky130_fd_sc_hd__a221o_1 _07255_ (.A1(net1268),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[20] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ),
    .C1(net1236),
    .X(_02685_));
 sky130_fd_sc_hd__o22a_1 _07256_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[20] ),
    .A2(net1219),
    .B1(_02684_),
    .B2(_02685_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__and3_1 _07257_ (.A(net1350),
    .B(net1363),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ),
    .X(_02686_));
 sky130_fd_sc_hd__a221o_1 _07258_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[21] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[21] ),
    .C1(net1237),
    .X(_02687_));
 sky130_fd_sc_hd__o22a_1 _07259_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[21] ),
    .A2(net1219),
    .B1(_02686_),
    .B2(_02687_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__and3_1 _07260_ (.A(net1348),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ),
    .X(_02688_));
 sky130_fd_sc_hd__a221o_1 _07261_ (.A1(net1270),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[22] ),
    .B1(net1155),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[22] ),
    .C1(net1237),
    .X(_02689_));
 sky130_fd_sc_hd__o22a_1 _07262_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[22] ),
    .A2(net1217),
    .B1(_02688_),
    .B2(_02689_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__and3_1 _07263_ (.A(net1348),
    .B(net1256),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[23] ),
    .X(_02690_));
 sky130_fd_sc_hd__a221o_1 _07264_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[23] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ),
    .C1(net1236),
    .X(_02691_));
 sky130_fd_sc_hd__o22a_1 _07265_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[23] ),
    .A2(net1218),
    .B1(_02690_),
    .B2(_02691_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__and3_1 _07266_ (.A(net1348),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ),
    .X(_02692_));
 sky130_fd_sc_hd__a221o_1 _07267_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[24] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[24] ),
    .C1(net1234),
    .X(_02693_));
 sky130_fd_sc_hd__o22a_1 _07268_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[24] ),
    .A2(net1217),
    .B1(_02692_),
    .B2(_02693_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__nor2_1 _07269_ (.A(_00958_),
    .B(net1211),
    .Y(_02694_));
 sky130_fd_sc_hd__a221o_1 _07270_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[25] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[25] ),
    .C1(net1234),
    .X(_02695_));
 sky130_fd_sc_hd__o22a_1 _07271_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[25] ),
    .A2(net1217),
    .B1(_02694_),
    .B2(_02695_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__nor2_1 _07272_ (.A(_00957_),
    .B(net1211),
    .Y(_02696_));
 sky130_fd_sc_hd__a221o_1 _07273_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[26] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[26] ),
    .C1(net1234),
    .X(_02697_));
 sky130_fd_sc_hd__o22a_1 _07274_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[26] ),
    .A2(net1217),
    .B1(_02696_),
    .B2(_02697_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__and3_1 _07275_ (.A(net1348),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ),
    .X(_02698_));
 sky130_fd_sc_hd__a221o_1 _07276_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[27] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[27] ),
    .C1(net1234),
    .X(_02699_));
 sky130_fd_sc_hd__o22a_1 _07277_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[27] ),
    .A2(net1217),
    .B1(_02698_),
    .B2(_02699_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__and3_1 _07278_ (.A(net1348),
    .B(net1362),
    .C(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ),
    .X(_02700_));
 sky130_fd_sc_hd__a221o_1 _07279_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[28] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[28] ),
    .C1(net1234),
    .X(_02701_));
 sky130_fd_sc_hd__o22a_1 _07280_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[28] ),
    .A2(net1217),
    .B1(_02700_),
    .B2(_02701_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__nor2_1 _07281_ (.A(_00956_),
    .B(net1211),
    .Y(_02702_));
 sky130_fd_sc_hd__a221o_1 _07282_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[29] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[29] ),
    .C1(net1234),
    .X(_02703_));
 sky130_fd_sc_hd__o22a_1 _07283_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[29] ),
    .A2(net1217),
    .B1(_02702_),
    .B2(_02703_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__nor2_1 _07284_ (.A(_00955_),
    .B(net1211),
    .Y(_02704_));
 sky130_fd_sc_hd__a221o_1 _07285_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[30] ),
    .B1(net1154),
    .B2(\u_pwm.u_pwm_2.u_reg.reg_2[30] ),
    .C1(net1234),
    .X(_02705_));
 sky130_fd_sc_hd__o22a_1 _07286_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[30] ),
    .A2(net1217),
    .B1(_02704_),
    .B2(_02705_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__and3_1 _07287_ (.A(net1348),
    .B(net1257),
    .C(\u_pwm.u_pwm_2.u_reg.reg_2[31] ),
    .X(_02706_));
 sky130_fd_sc_hd__a221o_1 _07288_ (.A1(net1266),
    .A2(\u_pwm.u_pwm_2.u_reg.reg_1[31] ),
    .B1(net1142),
    .B2(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ),
    .C1(net1234),
    .X(_02707_));
 sky130_fd_sc_hd__o22a_1 _07289_ (.A1(\u_pwm.u_pwm_2.u_reg.reg_0[31] ),
    .A2(net1217),
    .B1(_02706_),
    .B2(_02707_),
    .X(\u_pwm.u_pwm_2.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__and3_1 _07290_ (.A(net1355),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ),
    .X(_02708_));
 sky130_fd_sc_hd__a221o_1 _07291_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[0] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[0] ),
    .C1(net1240),
    .X(_02709_));
 sky130_fd_sc_hd__o22a_1 _07292_ (.A1(net2125),
    .A2(net1223),
    .B1(_02708_),
    .B2(_02709_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__and3_1 _07293_ (.A(net1355),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ),
    .X(_02710_));
 sky130_fd_sc_hd__a221o_1 _07294_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[1] ),
    .B1(net1158),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[1] ),
    .C1(net1239),
    .X(_02711_));
 sky130_fd_sc_hd__o22a_1 _07295_ (.A1(net2128),
    .A2(net1223),
    .B1(_02710_),
    .B2(_02711_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__and3_1 _07296_ (.A(net1355),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ),
    .X(_02712_));
 sky130_fd_sc_hd__a221o_1 _07297_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[2] ),
    .B1(net1157),
    .B2(net2101),
    .C1(net1240),
    .X(_02713_));
 sky130_fd_sc_hd__o22a_1 _07298_ (.A1(net2134),
    .A2(net1223),
    .B1(_02712_),
    .B2(_02713_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__nor2_1 _07299_ (.A(_00959_),
    .B(net1212),
    .Y(_02714_));
 sky130_fd_sc_hd__a221o_1 _07300_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[3] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[3] ),
    .C1(net1241),
    .X(_02715_));
 sky130_fd_sc_hd__o22a_1 _07301_ (.A1(net2123),
    .A2(net1224),
    .B1(_02714_),
    .B2(_02715_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__nor2_1 _07302_ (.A(_00960_),
    .B(net1212),
    .Y(_02716_));
 sky130_fd_sc_hd__a221o_1 _07303_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[4] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[4] ),
    .C1(net1240),
    .X(_02717_));
 sky130_fd_sc_hd__o22a_1 _07304_ (.A1(net2153),
    .A2(net1224),
    .B1(_02716_),
    .B2(_02717_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__and3_1 _07305_ (.A(net1355),
    .B(net1259),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[5] ),
    .X(_02718_));
 sky130_fd_sc_hd__a221o_1 _07306_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[5] ),
    .B1(net1143),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ),
    .C1(net1241),
    .X(_02719_));
 sky130_fd_sc_hd__o22a_1 _07307_ (.A1(net2077),
    .A2(net1224),
    .B1(_02718_),
    .B2(_02719_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__and3_1 _07308_ (.A(net1355),
    .B(net1258),
    .C(net2100),
    .X(_02720_));
 sky130_fd_sc_hd__a221o_1 _07309_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[6] ),
    .B1(net1143),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ),
    .C1(net1240),
    .X(_02721_));
 sky130_fd_sc_hd__o22a_1 _07310_ (.A1(net2103),
    .A2(net1223),
    .B1(_02720_),
    .B2(_02721_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__and3_1 _07311_ (.A(net1355),
    .B(net1258),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[7] ),
    .X(_02722_));
 sky130_fd_sc_hd__a221o_1 _07312_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[7] ),
    .B1(net1143),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ),
    .C1(net1240),
    .X(_02723_));
 sky130_fd_sc_hd__o22a_1 _07313_ (.A1(net2137),
    .A2(net1223),
    .B1(_02722_),
    .B2(_02723_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__nor2_1 _07314_ (.A(_00961_),
    .B(net1212),
    .Y(_02724_));
 sky130_fd_sc_hd__a221o_1 _07315_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[8] ),
    .B1(net1158),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[8] ),
    .C1(net1239),
    .X(_02725_));
 sky130_fd_sc_hd__o22a_1 _07316_ (.A1(net2183),
    .A2(net1223),
    .B1(_02724_),
    .B2(_02725_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__and3_1 _07317_ (.A(net1355),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ),
    .X(_02726_));
 sky130_fd_sc_hd__a221o_1 _07318_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[9] ),
    .B1(net1158),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[9] ),
    .C1(net1239),
    .X(_02727_));
 sky130_fd_sc_hd__o22a_1 _07319_ (.A1(net2147),
    .A2(net1223),
    .B1(_02726_),
    .B2(_02727_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__nor2_1 _07320_ (.A(_00962_),
    .B(net1213),
    .Y(_02728_));
 sky130_fd_sc_hd__a221o_1 _07321_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[10] ),
    .B1(net1158),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[10] ),
    .C1(net1239),
    .X(_02729_));
 sky130_fd_sc_hd__o22a_1 _07322_ (.A1(net2201),
    .A2(net1223),
    .B1(_02728_),
    .B2(_02729_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__nor2_1 _07323_ (.A(_00963_),
    .B(net1212),
    .Y(_02730_));
 sky130_fd_sc_hd__a221o_1 _07324_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[11] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[11] ),
    .C1(net1239),
    .X(_02731_));
 sky130_fd_sc_hd__o22a_1 _07325_ (.A1(net2140),
    .A2(net1223),
    .B1(_02730_),
    .B2(_02731_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__and3_1 _07326_ (.A(net1352),
    .B(net1372),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ),
    .X(_02732_));
 sky130_fd_sc_hd__a221o_1 _07327_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[12] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[12] ),
    .C1(net1241),
    .X(_02733_));
 sky130_fd_sc_hd__o22a_1 _07328_ (.A1(net2172),
    .A2(net1224),
    .B1(_02732_),
    .B2(_02733_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__and3_1 _07329_ (.A(net1352),
    .B(net1259),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[13] ),
    .X(_02734_));
 sky130_fd_sc_hd__a221o_1 _07330_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[13] ),
    .B1(net1143),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ),
    .C1(net1241),
    .X(_02735_));
 sky130_fd_sc_hd__o22a_1 _07331_ (.A1(net2217),
    .A2(net1224),
    .B1(_02734_),
    .B2(_02735_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__nor2_1 _07332_ (.A(_00965_),
    .B(net1212),
    .Y(_02736_));
 sky130_fd_sc_hd__a221o_1 _07333_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[14] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[14] ),
    .C1(net1241),
    .X(_02737_));
 sky130_fd_sc_hd__o22a_1 _07334_ (.A1(net2181),
    .A2(net1224),
    .B1(_02736_),
    .B2(_02737_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__and3_1 _07335_ (.A(net1352),
    .B(net1259),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[15] ),
    .X(_02738_));
 sky130_fd_sc_hd__a221o_1 _07336_ (.A1(net1273),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[15] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[15] ),
    .C1(net1239),
    .X(_02739_));
 sky130_fd_sc_hd__o22a_1 _07337_ (.A1(\u_pwm.u_pwm_1.u_reg.reg_0[15] ),
    .A2(net1223),
    .B1(_02738_),
    .B2(_02739_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__and3_1 _07338_ (.A(net1352),
    .B(net1363),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ),
    .X(_02740_));
 sky130_fd_sc_hd__a221o_1 _07339_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[16] ),
    .B1(net1156),
    .B2(net1974),
    .C1(net1237),
    .X(_02741_));
 sky130_fd_sc_hd__o22a_1 _07340_ (.A1(net2124),
    .A2(net1220),
    .B1(_02740_),
    .B2(_02741_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__and3_1 _07341_ (.A(net1352),
    .B(net1363),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .X(_02742_));
 sky130_fd_sc_hd__a221o_1 _07342_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[17] ),
    .B1(net1156),
    .B2(net1989),
    .C1(net1237),
    .X(_02743_));
 sky130_fd_sc_hd__o22a_1 _07343_ (.A1(net2194),
    .A2(net1220),
    .B1(_02742_),
    .B2(_02743_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__and3_1 _07344_ (.A(net1351),
    .B(net1256),
    .C(net1975),
    .X(_02744_));
 sky130_fd_sc_hd__a221o_1 _07345_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[18] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .C1(net1241),
    .X(_02745_));
 sky130_fd_sc_hd__o22a_1 _07346_ (.A1(net2204),
    .A2(net1224),
    .B1(_02744_),
    .B2(_02745_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__and3_1 _07347_ (.A(net1352),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .X(_02746_));
 sky130_fd_sc_hd__a221o_1 _07348_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[19] ),
    .B1(net1156),
    .B2(net1964),
    .C1(net1237),
    .X(_02747_));
 sky130_fd_sc_hd__o22a_1 _07349_ (.A1(net2092),
    .A2(net1220),
    .B1(_02746_),
    .B2(_02747_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__and3_1 _07350_ (.A(net1351),
    .B(net1256),
    .C(net1971),
    .X(_02748_));
 sky130_fd_sc_hd__a221o_1 _07351_ (.A1(net1274),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[20] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .C1(net1241),
    .X(_02749_));
 sky130_fd_sc_hd__o22a_1 _07352_ (.A1(net2226),
    .A2(net1224),
    .B1(_02748_),
    .B2(_02749_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__and3_1 _07353_ (.A(net1353),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ),
    .X(_02750_));
 sky130_fd_sc_hd__a221o_1 _07354_ (.A1(net1269),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[21] ),
    .B1(net1155),
    .B2(net1973),
    .C1(net1237),
    .X(_02751_));
 sky130_fd_sc_hd__o22a_1 _07355_ (.A1(net2156),
    .A2(net1220),
    .B1(_02750_),
    .B2(_02751_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__and3_1 _07356_ (.A(net1353),
    .B(net1364),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ),
    .X(_02752_));
 sky130_fd_sc_hd__a221o_1 _07357_ (.A1(net1270),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[22] ),
    .B1(net1156),
    .B2(net1972),
    .C1(net1237),
    .X(_02753_));
 sky130_fd_sc_hd__o22a_1 _07358_ (.A1(net2133),
    .A2(net1221),
    .B1(_02752_),
    .B2(_02753_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__and3_1 _07359_ (.A(net1351),
    .B(net1257),
    .C(net1987),
    .X(_02754_));
 sky130_fd_sc_hd__a221o_1 _07360_ (.A1(net1270),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[23] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ),
    .C1(net1237),
    .X(_02755_));
 sky130_fd_sc_hd__o22a_1 _07361_ (.A1(net2167),
    .A2(net1220),
    .B1(_02754_),
    .B2(_02755_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__and3_1 _07362_ (.A(net1352),
    .B(net1257),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[24] ),
    .X(_02756_));
 sky130_fd_sc_hd__a221o_1 _07363_ (.A1(net1271),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[24] ),
    .B1(net1143),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ),
    .C1(net1241),
    .X(_02757_));
 sky130_fd_sc_hd__o22a_1 _07364_ (.A1(net2188),
    .A2(net1222),
    .B1(_02756_),
    .B2(_02757_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__and3_1 _07365_ (.A(net1352),
    .B(net1363),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .X(_02758_));
 sky130_fd_sc_hd__a221o_1 _07366_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[25] ),
    .B1(net1159),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[25] ),
    .C1(net1235),
    .X(_02759_));
 sky130_fd_sc_hd__o22a_1 _07367_ (.A1(net2120),
    .A2(net1218),
    .B1(_02758_),
    .B2(_02759_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__and3_1 _07368_ (.A(net1352),
    .B(net1363),
    .C(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .X(_02760_));
 sky130_fd_sc_hd__a221o_1 _07369_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[26] ),
    .B1(net1156),
    .B2(net2127),
    .C1(net1235),
    .X(_02761_));
 sky130_fd_sc_hd__o22a_1 _07370_ (.A1(net2171),
    .A2(net1221),
    .B1(_02760_),
    .B2(_02761_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__nor2_1 _07371_ (.A(_00967_),
    .B(net1211),
    .Y(_02762_));
 sky130_fd_sc_hd__a221o_1 _07372_ (.A1(net1267),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[27] ),
    .B1(net1156),
    .B2(net2113),
    .C1(net1238),
    .X(_02763_));
 sky130_fd_sc_hd__o22a_1 _07373_ (.A1(net2192),
    .A2(net1221),
    .B1(_02762_),
    .B2(_02763_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__nor2_1 _07374_ (.A(_00968_),
    .B(net1211),
    .Y(_02764_));
 sky130_fd_sc_hd__a221o_1 _07375_ (.A1(net1271),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[28] ),
    .B1(net1156),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[28] ),
    .C1(net1237),
    .X(_02765_));
 sky130_fd_sc_hd__o22a_1 _07376_ (.A1(net2202),
    .A2(net1221),
    .B1(_02764_),
    .B2(_02765_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__nor2_1 _07377_ (.A(_00969_),
    .B(net1213),
    .Y(_02766_));
 sky130_fd_sc_hd__a221o_1 _07378_ (.A1(net1271),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[29] ),
    .B1(net1157),
    .B2(net2105),
    .C1(net1242),
    .X(_02767_));
 sky130_fd_sc_hd__o22a_1 _07379_ (.A1(net2158),
    .A2(net1222),
    .B1(_02766_),
    .B2(_02767_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__nor2_1 _07380_ (.A(_00970_),
    .B(net1213),
    .Y(_02768_));
 sky130_fd_sc_hd__a221o_1 _07381_ (.A1(net1271),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[30] ),
    .B1(net1157),
    .B2(\u_pwm.u_pwm_1.u_reg.reg_2[30] ),
    .C1(net1241),
    .X(_02769_));
 sky130_fd_sc_hd__o22a_1 _07382_ (.A1(net2214),
    .A2(net1222),
    .B1(_02768_),
    .B2(_02769_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__and3_1 _07383_ (.A(net1352),
    .B(net1259),
    .C(\u_pwm.u_pwm_1.u_reg.reg_2[31] ),
    .X(_02770_));
 sky130_fd_sc_hd__a221o_1 _07384_ (.A1(net1271),
    .A2(\u_pwm.u_pwm_1.u_reg.reg_1[31] ),
    .B1(net1144),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ),
    .C1(net1241),
    .X(_02771_));
 sky130_fd_sc_hd__o22a_1 _07385_ (.A1(net2191),
    .A2(net1222),
    .B1(_02770_),
    .B2(_02771_),
    .X(\u_pwm.u_pwm_1.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__xnor2_4 _07386_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .Y(_02772_));
 sky130_fd_sc_hd__xnor2_4 _07387_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .Y(_02773_));
 sky130_fd_sc_hd__or2_1 _07388_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ),
    .B(_02773_),
    .X(_02774_));
 sky130_fd_sc_hd__xnor2_4 _07389_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .Y(_02775_));
 sky130_fd_sc_hd__xnor2_2 _07390_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .Y(_02776_));
 sky130_fd_sc_hd__o211a_1 _07391_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ),
    .A2(_02775_),
    .B1(_02776_),
    .C1(\u_pwm.u_pwm_0.cfg_pwm_comp2[0] ),
    .X(_02777_));
 sky130_fd_sc_hd__xnor2_4 _07392_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ),
    .Y(_02778_));
 sky130_fd_sc_hd__a22o_1 _07393_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ),
    .A2(_02775_),
    .B1(_02778_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ),
    .X(_02779_));
 sky130_fd_sc_hd__xnor2_4 _07394_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ),
    .Y(_02780_));
 sky130_fd_sc_hd__or2_1 _07395_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ),
    .B(_02778_),
    .X(_02781_));
 sky130_fd_sc_hd__o221a_1 _07396_ (.A1(_02777_),
    .A2(_02779_),
    .B1(_02780_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ),
    .C1(_02781_),
    .X(_02782_));
 sky130_fd_sc_hd__xnor2_4 _07397_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .Y(_02783_));
 sky130_fd_sc_hd__a22o_1 _07398_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ),
    .A2(_02780_),
    .B1(_02783_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ),
    .X(_02784_));
 sky130_fd_sc_hd__xnor2_4 _07399_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ),
    .Y(_02785_));
 sky130_fd_sc_hd__o22a_1 _07400_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ),
    .A2(_02783_),
    .B1(_02785_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ),
    .X(_02786_));
 sky130_fd_sc_hd__o21a_1 _07401_ (.A1(_02782_),
    .A2(_02784_),
    .B1(_02786_),
    .X(_02787_));
 sky130_fd_sc_hd__xnor2_4 _07402_ (.A(net1077),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ),
    .Y(_02788_));
 sky130_fd_sc_hd__a22o_1 _07403_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ),
    .A2(_02785_),
    .B1(_02788_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ),
    .X(_02789_));
 sky130_fd_sc_hd__xnor2_4 _07404_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .Y(_02790_));
 sky130_fd_sc_hd__o22a_1 _07405_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ),
    .A2(_02788_),
    .B1(_02790_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ),
    .X(_02791_));
 sky130_fd_sc_hd__o21a_1 _07406_ (.A1(_02787_),
    .A2(_02789_),
    .B1(_02791_),
    .X(_02792_));
 sky130_fd_sc_hd__xnor2_4 _07407_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ),
    .Y(_02793_));
 sky130_fd_sc_hd__a221o_1 _07408_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ),
    .A2(_02790_),
    .B1(_02793_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ),
    .C1(_02792_),
    .X(_02794_));
 sky130_fd_sc_hd__xnor2_4 _07409_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .Y(_02795_));
 sky130_fd_sc_hd__o221a_1 _07410_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ),
    .A2(_02793_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ),
    .C1(_02794_),
    .X(_02796_));
 sky130_fd_sc_hd__a22o_1 _07411_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ),
    .A2(_02772_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ),
    .X(_02797_));
 sky130_fd_sc_hd__o221a_1 _07412_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ),
    .A2(_02772_),
    .B1(_02796_),
    .B2(_02797_),
    .C1(_02774_),
    .X(_02798_));
 sky130_fd_sc_hd__xnor2_4 _07413_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .Y(_02799_));
 sky130_fd_sc_hd__and2_1 _07414_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[14] ),
    .B(_02799_),
    .X(_02800_));
 sky130_fd_sc_hd__or2_1 _07415_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[14] ),
    .B(_02799_),
    .X(_02801_));
 sky130_fd_sc_hd__or3b_1 _07416_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ),
    .B(_02800_),
    .C_N(_02801_),
    .X(_02802_));
 sky130_fd_sc_hd__xnor2_4 _07417_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .Y(_02803_));
 sky130_fd_sc_hd__xnor2_4 _07418_ (.A(net1076),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .Y(_02804_));
 sky130_fd_sc_hd__o22ai_1 _07419_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ),
    .A2(_02803_),
    .B1(_02804_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ),
    .Y(_02805_));
 sky130_fd_sc_hd__and2_1 _07420_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ),
    .B(_02804_),
    .X(_02806_));
 sky130_fd_sc_hd__a221o_1 _07421_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ),
    .A2(_02773_),
    .B1(_02803_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ),
    .C1(_02806_),
    .X(_02807_));
 sky130_fd_sc_hd__or4_1 _07422_ (.A(_02798_),
    .B(_02802_),
    .C(_02805_),
    .D(_02807_),
    .X(_02808_));
 sky130_fd_sc_hd__nor2_1 _07423_ (.A(_02802_),
    .B(_02806_),
    .Y(_02809_));
 sky130_fd_sc_hd__o2bb2a_1 _07424_ (.A1_N(_02809_),
    .A2_N(_02805_),
    .B1(_02801_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ),
    .X(_02810_));
 sky130_fd_sc_hd__and2_1 _07425_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ),
    .X(_02811_));
 sky130_fd_sc_hd__and2_1 _07426_ (.A(_00860_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ),
    .X(_02812_));
 sky130_fd_sc_hd__nor2_1 _07427_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .B(_00940_),
    .Y(_02813_));
 sky130_fd_sc_hd__or2_1 _07428_ (.A(_02812_),
    .B(_02813_),
    .X(_02814_));
 sky130_fd_sc_hd__o22a_1 _07429_ (.A1(_00861_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ),
    .B2(_00860_),
    .X(_02815_));
 sky130_fd_sc_hd__a22o_1 _07430_ (.A1(_00862_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ),
    .B2(_00861_),
    .X(_02816_));
 sky130_fd_sc_hd__o22ai_1 _07431_ (.A1(_00863_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ),
    .B2(_00862_),
    .Y(_02817_));
 sky130_fd_sc_hd__a22o_1 _07432_ (.A1(_00864_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ),
    .B2(_00863_),
    .X(_02818_));
 sky130_fd_sc_hd__o22ai_1 _07433_ (.A1(_00865_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ),
    .B2(_00864_),
    .Y(_02819_));
 sky130_fd_sc_hd__and2b_1 _07434_ (.A_N(_02818_),
    .B(_02819_),
    .X(_02820_));
 sky130_fd_sc_hd__nor2_1 _07435_ (.A(_02817_),
    .B(_02820_),
    .Y(_02821_));
 sky130_fd_sc_hd__o21a_1 _07436_ (.A1(_02816_),
    .A2(_02821_),
    .B1(_02815_),
    .X(_02822_));
 sky130_fd_sc_hd__o211a_1 _07437_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[0] ),
    .C1(_00873_),
    .X(_02823_));
 sky130_fd_sc_hd__a221o_1 _07438_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ),
    .B2(_00871_),
    .C1(_02823_),
    .X(_02824_));
 sky130_fd_sc_hd__o221a_1 _07439_ (.A1(_00871_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ),
    .B2(_00870_),
    .C1(_02824_),
    .X(_02825_));
 sky130_fd_sc_hd__a221o_1 _07440_ (.A1(_00870_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ),
    .B2(_00869_),
    .C1(_02825_),
    .X(_02826_));
 sky130_fd_sc_hd__a22o_1 _07441_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ),
    .B2(net728),
    .X(_02827_));
 sky130_fd_sc_hd__o22a_1 _07442_ (.A1(_00869_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ),
    .B2(_00868_),
    .X(_02828_));
 sky130_fd_sc_hd__a21o_1 _07443_ (.A1(_02826_),
    .A2(_02828_),
    .B1(_02827_),
    .X(_02829_));
 sky130_fd_sc_hd__o221a_1 _07444_ (.A1(net728),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ),
    .B2(_00866_),
    .C1(_02829_),
    .X(_02830_));
 sky130_fd_sc_hd__a22o_1 _07445_ (.A1(_00866_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ),
    .B2(_00865_),
    .X(_02831_));
 sky130_fd_sc_hd__or2_1 _07446_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ),
    .X(_02832_));
 sky130_fd_sc_hd__or4_1 _07447_ (.A(_02816_),
    .B(_02817_),
    .C(_02818_),
    .D(_02819_),
    .X(_02833_));
 sky130_fd_sc_hd__a211o_1 _07448_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .A2(_00940_),
    .B1(_02811_),
    .C1(_02831_),
    .X(_02834_));
 sky130_fd_sc_hd__or4b_1 _07449_ (.A(_02812_),
    .B(_02834_),
    .C(_02813_),
    .D_N(_02815_),
    .X(_02835_));
 sky130_fd_sc_hd__or3_1 _07450_ (.A(_02830_),
    .B(_02833_),
    .C(_02835_),
    .X(_02836_));
 sky130_fd_sc_hd__o22a_1 _07451_ (.A1(_00859_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp2[14] ),
    .B1(_02814_),
    .B2(_02822_),
    .X(_02837_));
 sky130_fd_sc_hd__o2111a_1 _07452_ (.A1(_02811_),
    .A2(_02837_),
    .B1(_02832_),
    .C1(_00978_),
    .D1(_02836_),
    .X(_02838_));
 sky130_fd_sc_hd__a31o_1 _07453_ (.A1(\u_pwm.u_pwm_0.cfg_comp2_center ),
    .A2(_02808_),
    .A3(_02810_),
    .B1(_02838_),
    .X(_02839_));
 sky130_fd_sc_hd__o22a_1 _07454_ (.A1(_00858_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[15] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[14] ),
    .B2(_00859_),
    .X(_02840_));
 sky130_fd_sc_hd__nand2_1 _07455_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp0[15] ),
    .Y(_02841_));
 sky130_fd_sc_hd__and2b_1 _07456_ (.A_N(_02840_),
    .B(_02841_),
    .X(_02842_));
 sky130_fd_sc_hd__nand2_1 _07457_ (.A(_00860_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp0[13] ),
    .Y(_02843_));
 sky130_fd_sc_hd__o211a_1 _07458_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .A2(_00971_),
    .B1(_02840_),
    .C1(_02841_),
    .X(_02844_));
 sky130_fd_sc_hd__o22a_1 _07459_ (.A1(_00860_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[13] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ),
    .B2(_00861_),
    .X(_02845_));
 sky130_fd_sc_hd__inv_2 _07460_ (.A(_02845_),
    .Y(_02846_));
 sky130_fd_sc_hd__o22a_1 _07461_ (.A1(_00864_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ),
    .B2(_00865_),
    .X(_02847_));
 sky130_fd_sc_hd__o211a_1 _07462_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[0] ),
    .C1(_00873_),
    .X(_02848_));
 sky130_fd_sc_hd__a22o_1 _07463_ (.A1(_00871_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[2] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[1] ),
    .B2(_00872_),
    .X(_02849_));
 sky130_fd_sc_hd__o22a_1 _07464_ (.A1(_00870_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[3] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[2] ),
    .B2(_00871_),
    .X(_02850_));
 sky130_fd_sc_hd__o21a_1 _07465_ (.A1(_02848_),
    .A2(_02849_),
    .B1(_02850_),
    .X(_02851_));
 sky130_fd_sc_hd__a22o_1 _07466_ (.A1(_00869_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[4] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[3] ),
    .B2(_00870_),
    .X(_02852_));
 sky130_fd_sc_hd__o22a_1 _07467_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[5] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[4] ),
    .B2(_00869_),
    .X(_02853_));
 sky130_fd_sc_hd__o21a_1 _07468_ (.A1(_02851_),
    .A2(_02852_),
    .B1(_02853_),
    .X(_02854_));
 sky130_fd_sc_hd__a22o_1 _07469_ (.A1(net728),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[6] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[5] ),
    .B2(_00868_),
    .X(_02855_));
 sky130_fd_sc_hd__o22a_1 _07470_ (.A1(_00866_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[6] ),
    .B2(net728),
    .X(_02856_));
 sky130_fd_sc_hd__o21a_1 _07471_ (.A1(_02854_),
    .A2(_02855_),
    .B1(_02856_),
    .X(_02857_));
 sky130_fd_sc_hd__a22o_1 _07472_ (.A1(_00865_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[7] ),
    .B2(_00866_),
    .X(_02858_));
 sky130_fd_sc_hd__o21a_1 _07473_ (.A1(_02857_),
    .A2(_02858_),
    .B1(_02847_),
    .X(_02859_));
 sky130_fd_sc_hd__a22o_1 _07474_ (.A1(_00863_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ),
    .B2(_00864_),
    .X(_02860_));
 sky130_fd_sc_hd__o22a_1 _07475_ (.A1(_00862_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ),
    .B2(_00863_),
    .X(_02861_));
 sky130_fd_sc_hd__o21ai_1 _07476_ (.A1(_02859_),
    .A2(_02860_),
    .B1(_02861_),
    .Y(_02862_));
 sky130_fd_sc_hd__or2_1 _07477_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp0[14] ),
    .B(_02799_),
    .X(_02863_));
 sky130_fd_sc_hd__a22o_1 _07478_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ),
    .A2(_02803_),
    .B1(_02804_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[13] ),
    .X(_02864_));
 sky130_fd_sc_hd__o22a_1 _07479_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ),
    .A2(_02772_),
    .B1(_02773_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ),
    .X(_02865_));
 sky130_fd_sc_hd__a22o_1 _07480_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ),
    .A2(_02772_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ),
    .X(_02866_));
 sky130_fd_sc_hd__o22a_1 _07481_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ),
    .A2(_02793_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ),
    .X(_02867_));
 sky130_fd_sc_hd__or2_1 _07482_ (.A(_02866_),
    .B(_02867_),
    .X(_02868_));
 sky130_fd_sc_hd__a22o_1 _07483_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ),
    .A2(_02773_),
    .B1(_02865_),
    .B2(_02868_),
    .X(_02869_));
 sky130_fd_sc_hd__o211a_1 _07484_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[1] ),
    .A2(_02775_),
    .B1(_02776_),
    .C1(\u_pwm.u_pwm_0.cfg_pwm_comp0[0] ),
    .X(_02870_));
 sky130_fd_sc_hd__a22o_1 _07485_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[1] ),
    .A2(_02775_),
    .B1(_02778_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[2] ),
    .X(_02871_));
 sky130_fd_sc_hd__o22a_1 _07486_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[2] ),
    .A2(_02778_),
    .B1(_02780_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[3] ),
    .X(_02872_));
 sky130_fd_sc_hd__o21a_1 _07487_ (.A1(_02870_),
    .A2(_02871_),
    .B1(_02872_),
    .X(_02873_));
 sky130_fd_sc_hd__a22o_1 _07488_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[3] ),
    .A2(_02780_),
    .B1(_02783_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[4] ),
    .X(_02874_));
 sky130_fd_sc_hd__o22a_1 _07489_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[4] ),
    .A2(_02783_),
    .B1(_02785_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[5] ),
    .X(_02875_));
 sky130_fd_sc_hd__o21a_1 _07490_ (.A1(_02873_),
    .A2(_02874_),
    .B1(_02875_),
    .X(_02876_));
 sky130_fd_sc_hd__a22o_1 _07491_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[5] ),
    .A2(_02785_),
    .B1(_02788_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[6] ),
    .X(_02877_));
 sky130_fd_sc_hd__or2_1 _07492_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp0[7] ),
    .B(_02790_),
    .X(_02878_));
 sky130_fd_sc_hd__o221a_1 _07493_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[6] ),
    .A2(_02788_),
    .B1(_02876_),
    .B2(_02877_),
    .C1(_02878_),
    .X(_02879_));
 sky130_fd_sc_hd__a22o_1 _07494_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ),
    .A2(_02773_),
    .B1(_02790_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[7] ),
    .X(_02880_));
 sky130_fd_sc_hd__a2bb2o_1 _07495_ (.A1_N(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ),
    .A2_N(_02803_),
    .B1(_02793_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ),
    .X(_02881_));
 sky130_fd_sc_hd__nand2_1 _07496_ (.A(_02865_),
    .B(_02867_),
    .Y(_02882_));
 sky130_fd_sc_hd__or4_1 _07497_ (.A(_02866_),
    .B(_02880_),
    .C(_02881_),
    .D(_02882_),
    .X(_02883_));
 sky130_fd_sc_hd__o221a_1 _07498_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ),
    .A2(_02803_),
    .B1(_02879_),
    .B2(_02883_),
    .C1(_02869_),
    .X(_02884_));
 sky130_fd_sc_hd__o221a_1 _07499_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[13] ),
    .A2(_02804_),
    .B1(_02864_),
    .B2(_02884_),
    .C1(_02863_),
    .X(_02885_));
 sky130_fd_sc_hd__o221a_1 _07500_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .A2(_00972_),
    .B1(_00973_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .C1(_02843_),
    .X(_02886_));
 sky130_fd_sc_hd__and4_1 _07501_ (.A(_02844_),
    .B(_02845_),
    .C(_02862_),
    .D(_02886_),
    .X(_02887_));
 sky130_fd_sc_hd__a311o_1 _07502_ (.A1(_02843_),
    .A2(_02844_),
    .A3(_02846_),
    .B1(_02842_),
    .C1(\u_pwm.u_pwm_0.cfg_comp0_center ),
    .X(_02888_));
 sky130_fd_sc_hd__a211o_1 _07503_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp0[14] ),
    .A2(_02799_),
    .B1(_02885_),
    .C1(\u_pwm.u_pwm_0.cfg_pwm_comp0[15] ),
    .X(_02889_));
 sky130_fd_sc_hd__o2bb2a_1 _07504_ (.A1_N(\u_pwm.u_pwm_0.cfg_comp0_center ),
    .A2_N(_02889_),
    .B1(_02888_),
    .B2(_02887_),
    .X(_02890_));
 sky130_fd_sc_hd__a2bb2o_1 _07505_ (.A1_N(_00862_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_comp1[11] ),
    .B1(_00975_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .X(_02891_));
 sky130_fd_sc_hd__nand2_1 _07506_ (.A(_00865_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp1[8] ),
    .Y(_02892_));
 sky130_fd_sc_hd__o211a_1 _07507_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[0] ),
    .C1(_00873_),
    .X(_02893_));
 sky130_fd_sc_hd__a22o_1 _07508_ (.A1(_00871_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[2] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[1] ),
    .B2(_00872_),
    .X(_02894_));
 sky130_fd_sc_hd__o22a_1 _07509_ (.A1(_00870_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[3] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[2] ),
    .B2(_00871_),
    .X(_02895_));
 sky130_fd_sc_hd__o21a_1 _07510_ (.A1(_02893_),
    .A2(_02894_),
    .B1(_02895_),
    .X(_02896_));
 sky130_fd_sc_hd__a22o_1 _07511_ (.A1(_00869_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[4] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[3] ),
    .B2(_00870_),
    .X(_02897_));
 sky130_fd_sc_hd__o22a_1 _07512_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[5] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[4] ),
    .B2(_00869_),
    .X(_02898_));
 sky130_fd_sc_hd__o21a_1 _07513_ (.A1(_02896_),
    .A2(_02897_),
    .B1(_02898_),
    .X(_02899_));
 sky130_fd_sc_hd__a22o_1 _07514_ (.A1(_00866_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[5] ),
    .B2(_00868_),
    .X(_02900_));
 sky130_fd_sc_hd__a21o_1 _07515_ (.A1(net728),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ),
    .B1(_02900_),
    .X(_02901_));
 sky130_fd_sc_hd__o22a_1 _07516_ (.A1(_00866_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ),
    .B2(net728),
    .X(_02902_));
 sky130_fd_sc_hd__o21ai_1 _07517_ (.A1(_02899_),
    .A2(_02901_),
    .B1(_02902_),
    .Y(_02903_));
 sky130_fd_sc_hd__or4_1 _07518_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .B(net728),
    .C(_00977_),
    .D(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ),
    .X(_02904_));
 sky130_fd_sc_hd__a2bb2o_1 _07519_ (.A1_N(\u_pwm.u_pwm_0.cfg_pwm_comp1[8] ),
    .A2_N(_00865_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .B2(_00976_),
    .X(_02905_));
 sky130_fd_sc_hd__a31o_1 _07520_ (.A1(_02892_),
    .A2(_02903_),
    .A3(_02904_),
    .B1(_02905_),
    .X(_02906_));
 sky130_fd_sc_hd__o221a_1 _07521_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .A2(_00975_),
    .B1(_00976_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .C1(_02906_),
    .X(_02907_));
 sky130_fd_sc_hd__o22a_1 _07522_ (.A1(_00858_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[15] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ),
    .B2(_00859_),
    .X(_02908_));
 sky130_fd_sc_hd__nand2_1 _07523_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp1[15] ),
    .Y(_02909_));
 sky130_fd_sc_hd__o211a_1 _07524_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .A2(_00974_),
    .B1(_02908_),
    .C1(_02909_),
    .X(_02910_));
 sky130_fd_sc_hd__o22ai_1 _07525_ (.A1(_00860_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[13] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp1[12] ),
    .B2(_00861_),
    .Y(_02911_));
 sky130_fd_sc_hd__nand2_1 _07526_ (.A(_00861_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp1[12] ),
    .Y(_02912_));
 sky130_fd_sc_hd__nand2_1 _07527_ (.A(_00860_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp1[13] ),
    .Y(_02913_));
 sky130_fd_sc_hd__nand2_1 _07528_ (.A(_00862_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp1[11] ),
    .Y(_02914_));
 sky130_fd_sc_hd__and3b_1 _07529_ (.A_N(_02911_),
    .B(_02912_),
    .C(_02913_),
    .X(_02915_));
 sky130_fd_sc_hd__o2111a_1 _07530_ (.A1(_02891_),
    .A2(_02907_),
    .B1(_02910_),
    .C1(_02914_),
    .D1(_02915_),
    .X(_02916_));
 sky130_fd_sc_hd__and2b_1 _07531_ (.A_N(_02908_),
    .B(_02909_),
    .X(_02917_));
 sky130_fd_sc_hd__o22a_1 _07532_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[12] ),
    .A2(_02803_),
    .B1(_02804_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[13] ),
    .X(_02918_));
 sky130_fd_sc_hd__a22oi_1 _07533_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[11] ),
    .A2(_02773_),
    .B1(_02803_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[12] ),
    .Y(_02919_));
 sky130_fd_sc_hd__o22a_1 _07534_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[10] ),
    .A2(_02772_),
    .B1(_02773_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[11] ),
    .X(_02920_));
 sky130_fd_sc_hd__a22o_1 _07535_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[10] ),
    .A2(_02772_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[9] ),
    .X(_02921_));
 sky130_fd_sc_hd__o22a_1 _07536_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[8] ),
    .A2(_02793_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[9] ),
    .X(_02922_));
 sky130_fd_sc_hd__o211a_1 _07537_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[1] ),
    .A2(_02775_),
    .B1(_02776_),
    .C1(\u_pwm.u_pwm_0.cfg_pwm_comp1[0] ),
    .X(_02923_));
 sky130_fd_sc_hd__a22o_1 _07538_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[1] ),
    .A2(_02775_),
    .B1(_02778_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[2] ),
    .X(_02924_));
 sky130_fd_sc_hd__or2_1 _07539_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[2] ),
    .B(_02778_),
    .X(_02925_));
 sky130_fd_sc_hd__o221a_1 _07540_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[3] ),
    .A2(_02780_),
    .B1(_02923_),
    .B2(_02924_),
    .C1(_02925_),
    .X(_02926_));
 sky130_fd_sc_hd__a22o_1 _07541_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[3] ),
    .A2(_02780_),
    .B1(_02783_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[4] ),
    .X(_02927_));
 sky130_fd_sc_hd__o22a_1 _07542_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[4] ),
    .A2(_02783_),
    .B1(_02785_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[5] ),
    .X(_02928_));
 sky130_fd_sc_hd__o21a_1 _07543_ (.A1(_02926_),
    .A2(_02927_),
    .B1(_02928_),
    .X(_02929_));
 sky130_fd_sc_hd__a221o_1 _07544_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[5] ),
    .A2(_02785_),
    .B1(_02788_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ),
    .C1(_02929_),
    .X(_02930_));
 sky130_fd_sc_hd__o22a_1 _07545_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ),
    .A2(_02788_),
    .B1(_02790_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ),
    .X(_02931_));
 sky130_fd_sc_hd__o21ai_1 _07546_ (.A1(_02921_),
    .A2(_02922_),
    .B1(_02920_),
    .Y(_02932_));
 sky130_fd_sc_hd__nand2_1 _07547_ (.A(_02919_),
    .B(_02932_),
    .Y(_02933_));
 sky130_fd_sc_hd__a221o_1 _07548_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ),
    .A2(_02790_),
    .B1(_02793_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[8] ),
    .C1(_02921_),
    .X(_02934_));
 sky130_fd_sc_hd__nand4_1 _07549_ (.A(_02918_),
    .B(_02919_),
    .C(_02920_),
    .D(_02922_),
    .Y(_02935_));
 sky130_fd_sc_hd__a211o_1 _07550_ (.A1(_02930_),
    .A2(_02931_),
    .B1(_02934_),
    .C1(_02935_),
    .X(_02936_));
 sky130_fd_sc_hd__nor2_1 _07551_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ),
    .B(_02799_),
    .Y(_02937_));
 sky130_fd_sc_hd__and2_1 _07552_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ),
    .B(_02799_),
    .X(_02938_));
 sky130_fd_sc_hd__a32o_1 _07553_ (.A1(_02918_),
    .A2(_02933_),
    .A3(_02936_),
    .B1(_02804_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp1[13] ),
    .X(_02939_));
 sky130_fd_sc_hd__or4_1 _07554_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp1[15] ),
    .B(_02937_),
    .C(_02938_),
    .D(_02939_),
    .X(_02940_));
 sky130_fd_sc_hd__o31a_1 _07555_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp1[15] ),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ),
    .A3(_02799_),
    .B1(\u_pwm.u_pwm_0.cfg_comp1_center ),
    .X(_02941_));
 sky130_fd_sc_hd__a311o_1 _07556_ (.A1(_02910_),
    .A2(_02911_),
    .A3(_02913_),
    .B1(_02917_),
    .C1(\u_pwm.u_pwm_0.cfg_comp1_center ),
    .X(_02942_));
 sky130_fd_sc_hd__a2bb2o_1 _07557_ (.A1_N(_02916_),
    .A2_N(_02942_),
    .B1(_02940_),
    .B2(_02941_),
    .X(_02943_));
 sky130_fd_sc_hd__xnor2_1 _07558_ (.A(_02890_),
    .B(_02943_),
    .Y(_02944_));
 sky130_fd_sc_hd__xor2_1 _07559_ (.A(_02839_),
    .B(_02944_),
    .X(_02945_));
 sky130_fd_sc_hd__and2_1 _07560_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ),
    .X(_02946_));
 sky130_fd_sc_hd__nor2_1 _07561_ (.A(_00859_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .Y(_02947_));
 sky130_fd_sc_hd__a22o_1 _07562_ (.A1(_00860_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .B2(_00859_),
    .X(_02948_));
 sky130_fd_sc_hd__o22ai_1 _07563_ (.A1(_00861_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ),
    .B2(_00860_),
    .Y(_02949_));
 sky130_fd_sc_hd__a2bb2o_1 _07564_ (.A1_N(_00862_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .B2(_00942_),
    .X(_02950_));
 sky130_fd_sc_hd__nand2_1 _07565_ (.A(_00861_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ),
    .Y(_02951_));
 sky130_fd_sc_hd__nand2_1 _07566_ (.A(_00862_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .Y(_02952_));
 sky130_fd_sc_hd__nand2_1 _07567_ (.A(_02951_),
    .B(_02952_),
    .Y(_02953_));
 sky130_fd_sc_hd__a2bb2o_1 _07568_ (.A1_N(_00865_),
    .A2_N(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ),
    .B1(_00941_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .X(_02954_));
 sky130_fd_sc_hd__o221a_1 _07569_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .A2(_00941_),
    .B1(_00942_),
    .B2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .C1(_02954_),
    .X(_02955_));
 sky130_fd_sc_hd__o211a_1 _07570_ (.A1(_02950_),
    .A2(_02955_),
    .B1(_02952_),
    .C1(_02951_),
    .X(_02956_));
 sky130_fd_sc_hd__nor2_1 _07571_ (.A(_02949_),
    .B(_02956_),
    .Y(_02957_));
 sky130_fd_sc_hd__o21ba_1 _07572_ (.A1(_02948_),
    .A2(_02957_),
    .B1_N(_02947_),
    .X(_02958_));
 sky130_fd_sc_hd__o211a_1 _07573_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ),
    .C1(_00873_),
    .X(_02959_));
 sky130_fd_sc_hd__a221o_1 _07574_ (.A1(_00872_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ),
    .B2(_00871_),
    .C1(_02959_),
    .X(_02960_));
 sky130_fd_sc_hd__o221a_1 _07575_ (.A1(_00871_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ),
    .B2(_00870_),
    .C1(_02960_),
    .X(_02961_));
 sky130_fd_sc_hd__a221o_1 _07576_ (.A1(_00870_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ),
    .B2(_00869_),
    .C1(_02961_),
    .X(_02962_));
 sky130_fd_sc_hd__o221a_1 _07577_ (.A1(_00869_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ),
    .B2(_00868_),
    .C1(_02962_),
    .X(_02963_));
 sky130_fd_sc_hd__a221o_1 _07578_ (.A1(_00868_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ),
    .B2(net728),
    .C1(_02963_),
    .X(_02964_));
 sky130_fd_sc_hd__o221a_1 _07579_ (.A1(_00867_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ),
    .B2(_00866_),
    .C1(_02964_),
    .X(_02965_));
 sky130_fd_sc_hd__a221o_1 _07580_ (.A1(_00864_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[9] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ),
    .B2(_00863_),
    .C1(_02949_),
    .X(_02966_));
 sky130_fd_sc_hd__a221o_1 _07581_ (.A1(_00866_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ),
    .B2(_00865_),
    .C1(_02946_),
    .X(_02967_));
 sky130_fd_sc_hd__nor2_1 _07582_ (.A(_00858_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ),
    .Y(_02968_));
 sky130_fd_sc_hd__or4_1 _07583_ (.A(_02947_),
    .B(_02953_),
    .C(_02967_),
    .D(_02968_),
    .X(_02969_));
 sky130_fd_sc_hd__or3_1 _07584_ (.A(_02950_),
    .B(_02954_),
    .C(_02969_),
    .X(_02970_));
 sky130_fd_sc_hd__or4_1 _07585_ (.A(_02948_),
    .B(_02965_),
    .C(_02966_),
    .D(_02970_),
    .X(_02971_));
 sky130_fd_sc_hd__nor2_1 _07586_ (.A(\u_pwm.u_pwm_0.cfg_comp3_center ),
    .B(_02968_),
    .Y(_02972_));
 sky130_fd_sc_hd__o211a_1 _07587_ (.A1(_02946_),
    .A2(_02958_),
    .B1(_02971_),
    .C1(_02972_),
    .X(_02973_));
 sky130_fd_sc_hd__or2_1 _07588_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ),
    .B(_02803_),
    .X(_02974_));
 sky130_fd_sc_hd__and2_1 _07589_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ),
    .B(_02803_),
    .X(_02975_));
 sky130_fd_sc_hd__o22a_1 _07590_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ),
    .A2(_02772_),
    .B1(_02773_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .X(_02976_));
 sky130_fd_sc_hd__a22o_1 _07591_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ),
    .A2(_02772_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[9] ),
    .X(_02977_));
 sky130_fd_sc_hd__o22a_1 _07592_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ),
    .A2(_02793_),
    .B1(_02795_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[9] ),
    .X(_02978_));
 sky130_fd_sc_hd__nand2_1 _07593_ (.A(_02976_),
    .B(_02978_),
    .Y(_02979_));
 sky130_fd_sc_hd__or2_1 _07594_ (.A(_02977_),
    .B(_02978_),
    .X(_02980_));
 sky130_fd_sc_hd__a22o_1 _07595_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .A2(_02773_),
    .B1(_02976_),
    .B2(_02980_),
    .X(_02981_));
 sky130_fd_sc_hd__o211a_1 _07596_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ),
    .A2(_02775_),
    .B1(_02776_),
    .C1(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ),
    .X(_02982_));
 sky130_fd_sc_hd__a22o_1 _07597_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ),
    .A2(_02775_),
    .B1(_02778_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ),
    .X(_02983_));
 sky130_fd_sc_hd__o22a_1 _07598_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ),
    .A2(_02778_),
    .B1(_02780_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ),
    .X(_02984_));
 sky130_fd_sc_hd__o21a_1 _07599_ (.A1(_02982_),
    .A2(_02983_),
    .B1(_02984_),
    .X(_02985_));
 sky130_fd_sc_hd__a221o_1 _07600_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ),
    .A2(_02780_),
    .B1(_02783_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ),
    .C1(_02985_),
    .X(_02986_));
 sky130_fd_sc_hd__o221a_1 _07601_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ),
    .A2(_02783_),
    .B1(_02785_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ),
    .C1(_02986_),
    .X(_02987_));
 sky130_fd_sc_hd__a221o_1 _07602_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ),
    .A2(_02785_),
    .B1(_02788_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ),
    .C1(_02987_),
    .X(_02988_));
 sky130_fd_sc_hd__o221a_1 _07603_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ),
    .A2(_02788_),
    .B1(_02790_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ),
    .C1(_02988_),
    .X(_02989_));
 sky130_fd_sc_hd__a22o_1 _07604_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ),
    .A2(_02773_),
    .B1(_02790_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ),
    .X(_02990_));
 sky130_fd_sc_hd__a211o_1 _07605_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ),
    .A2(_02793_),
    .B1(_02977_),
    .C1(_02990_),
    .X(_02991_));
 sky130_fd_sc_hd__o31a_1 _07606_ (.A1(_02979_),
    .A2(_02989_),
    .A3(_02991_),
    .B1(_02981_),
    .X(_02992_));
 sky130_fd_sc_hd__o221a_1 _07607_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ),
    .A2(_02804_),
    .B1(_02975_),
    .B2(_02992_),
    .C1(_02974_),
    .X(_02993_));
 sky130_fd_sc_hd__nor2_1 _07608_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .B(_02799_),
    .Y(_02994_));
 sky130_fd_sc_hd__a22o_1 _07609_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .A2(_02799_),
    .B1(_02804_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ),
    .X(_02995_));
 sky130_fd_sc_hd__or4_1 _07610_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ),
    .B(_02993_),
    .C(_02994_),
    .D(_02995_),
    .X(_02996_));
 sky130_fd_sc_hd__or3_1 _07611_ (.A(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ),
    .C(_02799_),
    .X(_02997_));
 sky130_fd_sc_hd__a31o_1 _07612_ (.A1(\u_pwm.u_pwm_0.cfg_comp3_center ),
    .A2(_02996_),
    .A3(_02997_),
    .B1(_02973_),
    .X(_02998_));
 sky130_fd_sc_hd__nand2_1 _07613_ (.A(_02945_),
    .B(_02998_),
    .Y(_02999_));
 sky130_fd_sc_hd__or2_1 _07614_ (.A(_02945_),
    .B(_02998_),
    .X(_03000_));
 sky130_fd_sc_hd__and4_1 _07615_ (.A(\u_pwm.u_pwm_0.cfg_pwm_mode[1] ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_mode[0] ),
    .C(_02999_),
    .D(_03000_),
    .X(_03001_));
 sky130_fd_sc_hd__and2b_1 _07616_ (.A_N(_02944_),
    .B(\u_pwm.u_pwm_0.cfg_pwm_mode[0] ),
    .X(_03002_));
 sky130_fd_sc_hd__o22ai_1 _07617_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_mode[0] ),
    .A2(_02945_),
    .B1(_03002_),
    .B2(\u_pwm.u_pwm_0.cfg_pwm_mode[1] ),
    .Y(_03003_));
 sky130_fd_sc_hd__o32a_1 _07618_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_mode[1] ),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_mode[0] ),
    .A3(_02890_),
    .B1(_03001_),
    .B2(_03003_),
    .X(\u_pwm.u_pwm_0.u_pwm.pwm_wfm_i ));
 sky130_fd_sc_hd__xnor2_4 _07619_ (.A(net1075),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .Y(_03004_));
 sky130_fd_sc_hd__a21oi_2 _07620_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[14] ),
    .A2(_03004_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[15] ),
    .Y(_03005_));
 sky130_fd_sc_hd__xnor2_4 _07621_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ),
    .Y(_03006_));
 sky130_fd_sc_hd__xnor2_4 _07622_ (.A(net1075),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .Y(_03007_));
 sky130_fd_sc_hd__xnor2_4 _07623_ (.A(net1075),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .Y(_03008_));
 sky130_fd_sc_hd__a22o_1 _07624_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[13] ),
    .A2(_03007_),
    .B1(_03008_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[12] ),
    .X(_03009_));
 sky130_fd_sc_hd__xnor2_4 _07625_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .Y(_03010_));
 sky130_fd_sc_hd__xnor2_4 _07626_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .Y(_03011_));
 sky130_fd_sc_hd__o22a_1 _07627_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[9] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ),
    .X(_03012_));
 sky130_fd_sc_hd__and2b_1 _07628_ (.A_N(_03009_),
    .B(_03012_),
    .X(_03013_));
 sky130_fd_sc_hd__a22o_1 _07629_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ),
    .A2(_03006_),
    .B1(_03010_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[9] ),
    .X(_03014_));
 sky130_fd_sc_hd__xnor2_4 _07630_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .Y(_03015_));
 sky130_fd_sc_hd__a22o_1 _07631_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ),
    .A2(_03011_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[11] ),
    .X(_03016_));
 sky130_fd_sc_hd__o22a_1 _07632_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[12] ),
    .A2(_03008_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[11] ),
    .X(_03017_));
 sky130_fd_sc_hd__o22a_1 _07633_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[14] ),
    .A2(_03004_),
    .B1(_03007_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[13] ),
    .X(_03018_));
 sky130_fd_sc_hd__and4bb_1 _07634_ (.A_N(_03014_),
    .B_N(_03016_),
    .C(_03017_),
    .D(_03018_),
    .X(_03019_));
 sky130_fd_sc_hd__o2111ai_4 _07635_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ),
    .A2(_03006_),
    .B1(_03013_),
    .C1(_03019_),
    .D1(_03005_),
    .Y(_03020_));
 sky130_fd_sc_hd__xnor2_4 _07636_ (.A(net1075),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .Y(_03021_));
 sky130_fd_sc_hd__xnor2_4 _07637_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .Y(_03022_));
 sky130_fd_sc_hd__o22a_1 _07638_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ),
    .X(_03023_));
 sky130_fd_sc_hd__nand2_1 _07639_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ),
    .B(_03022_),
    .Y(_03024_));
 sky130_fd_sc_hd__and2b_1 _07640_ (.A_N(_03023_),
    .B(_03024_),
    .X(_03025_));
 sky130_fd_sc_hd__xnor2_4 _07641_ (.A(net1075),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ),
    .Y(_03026_));
 sky130_fd_sc_hd__xnor2_4 _07642_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ),
    .Y(_03027_));
 sky130_fd_sc_hd__a22o_1 _07643_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ),
    .A2(_03026_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ),
    .X(_03028_));
 sky130_fd_sc_hd__or2_1 _07644_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ),
    .B(_03027_),
    .X(_03029_));
 sky130_fd_sc_hd__xnor2_4 _07645_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .Y(_03030_));
 sky130_fd_sc_hd__xnor2_4 _07646_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[5] ),
    .Y(_03031_));
 sky130_fd_sc_hd__a22o_1 _07647_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[4] ),
    .A2(_03030_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ),
    .X(_03032_));
 sky130_fd_sc_hd__or2_1 _07648_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ),
    .B(_03031_),
    .X(_03033_));
 sky130_fd_sc_hd__or2_1 _07649_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ),
    .B(_03026_),
    .X(_03034_));
 sky130_fd_sc_hd__and4b_1 _07650_ (.A_N(_03028_),
    .B(_03029_),
    .C(_03033_),
    .D(_03034_),
    .X(_03035_));
 sky130_fd_sc_hd__o21ai_1 _07651_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[4] ),
    .A2(_03030_),
    .B1(_03035_),
    .Y(_03036_));
 sky130_fd_sc_hd__nor2_1 _07652_ (.A(_03032_),
    .B(_03036_),
    .Y(_03037_));
 sky130_fd_sc_hd__xnor2_1 _07653_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .Y(_03038_));
 sky130_fd_sc_hd__and2_1 _07654_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ),
    .B(net588),
    .X(_03039_));
 sky130_fd_sc_hd__nor2_1 _07655_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ),
    .B(net588),
    .Y(_03040_));
 sky130_fd_sc_hd__xnor2_1 _07656_ (.A(net1074),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .Y(_03041_));
 sky130_fd_sc_hd__and2_1 _07657_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ),
    .B(net587),
    .X(_03042_));
 sky130_fd_sc_hd__nor2_1 _07658_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ),
    .B(net587),
    .Y(_03043_));
 sky130_fd_sc_hd__or4_1 _07659_ (.A(_03039_),
    .B(_03040_),
    .C(_03042_),
    .D(_03043_),
    .X(_03044_));
 sky130_fd_sc_hd__o211a_1 _07660_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ),
    .A2(net587),
    .B1(net588),
    .C1(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ),
    .X(_03045_));
 sky130_fd_sc_hd__nor2_1 _07661_ (.A(_03025_),
    .B(_03044_),
    .Y(_03046_));
 sky130_fd_sc_hd__o31a_1 _07662_ (.A1(_03042_),
    .A2(_03045_),
    .A3(_03046_),
    .B1(_03037_),
    .X(_03047_));
 sky130_fd_sc_hd__a221oi_1 _07663_ (.A1(_03028_),
    .A2(_03029_),
    .B1(_03032_),
    .B2(_03035_),
    .C1(_03047_),
    .Y(_03048_));
 sky130_fd_sc_hd__a21o_1 _07664_ (.A1(_03012_),
    .A2(_03014_),
    .B1(_03016_),
    .X(_03049_));
 sky130_fd_sc_hd__a21o_1 _07665_ (.A1(_03017_),
    .A2(_03049_),
    .B1(_03009_),
    .X(_03050_));
 sky130_fd_sc_hd__nand2_1 _07666_ (.A(_03018_),
    .B(_03050_),
    .Y(_03051_));
 sky130_fd_sc_hd__o211a_1 _07667_ (.A1(_03020_),
    .A2(_03048_),
    .B1(_03051_),
    .C1(_03005_),
    .X(_03052_));
 sky130_fd_sc_hd__a211oi_1 _07668_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ),
    .A2(_03021_),
    .B1(_03044_),
    .C1(_03020_),
    .Y(_03053_));
 sky130_fd_sc_hd__a41o_1 _07669_ (.A1(_03023_),
    .A2(_03024_),
    .A3(_03037_),
    .A4(_03053_),
    .B1(_00981_),
    .X(_03054_));
 sky130_fd_sc_hd__a22o_1 _07670_ (.A1(net727),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[15] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[14] ),
    .B2(_00879_),
    .X(_03055_));
 sky130_fd_sc_hd__o22ai_1 _07671_ (.A1(net727),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[15] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[13] ),
    .B2(_00880_),
    .Y(_03056_));
 sky130_fd_sc_hd__a211o_1 _07672_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .A2(_00980_),
    .B1(_03055_),
    .C1(_03056_),
    .X(_03057_));
 sky130_fd_sc_hd__nand2_1 _07673_ (.A(_00882_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[11] ),
    .Y(_03058_));
 sky130_fd_sc_hd__nand2_1 _07674_ (.A(_00883_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ),
    .Y(_03059_));
 sky130_fd_sc_hd__nand2_1 _07675_ (.A(_03058_),
    .B(_03059_),
    .Y(_03060_));
 sky130_fd_sc_hd__or2_1 _07676_ (.A(_00882_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[11] ),
    .X(_03061_));
 sky130_fd_sc_hd__or2_1 _07677_ (.A(_00884_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[9] ),
    .X(_03062_));
 sky130_fd_sc_hd__o21a_1 _07678_ (.A1(_00883_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ),
    .B1(_03058_),
    .X(_03063_));
 sky130_fd_sc_hd__and3_1 _07679_ (.A(_03059_),
    .B(_03061_),
    .C(_03063_),
    .X(_03064_));
 sky130_fd_sc_hd__nand2_1 _07680_ (.A(_03062_),
    .B(_03064_),
    .Y(_03065_));
 sky130_fd_sc_hd__a22o_1 _07681_ (.A1(_00884_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[9] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ),
    .B2(_00885_),
    .X(_03066_));
 sky130_fd_sc_hd__a22o_1 _07682_ (.A1(_00880_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[13] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[12] ),
    .B2(_00881_),
    .X(_03067_));
 sky130_fd_sc_hd__or2_1 _07683_ (.A(_00881_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[12] ),
    .X(_03068_));
 sky130_fd_sc_hd__nor2_1 _07684_ (.A(_00885_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ),
    .Y(_03069_));
 sky130_fd_sc_hd__or3b_1 _07685_ (.A(_03069_),
    .B(_03067_),
    .C_N(_03068_),
    .X(_03070_));
 sky130_fd_sc_hd__or4_1 _07686_ (.A(_03057_),
    .B(_03065_),
    .C(_03066_),
    .D(_03070_),
    .X(_03071_));
 sky130_fd_sc_hd__a22o_1 _07687_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp0[4] ),
    .B2(_00889_),
    .X(_03072_));
 sky130_fd_sc_hd__nor2_1 _07688_ (.A(_00889_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[4] ),
    .Y(_03073_));
 sky130_fd_sc_hd__nand2b_1 _07689_ (.A_N(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ),
    .Y(_03074_));
 sky130_fd_sc_hd__nand2b_1 _07690_ (.A_N(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .Y(_03075_));
 sky130_fd_sc_hd__xnor2_1 _07691_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ),
    .Y(_03076_));
 sky130_fd_sc_hd__and3_1 _07692_ (.A(_03074_),
    .B(_03075_),
    .C(_03076_),
    .X(_03077_));
 sky130_fd_sc_hd__a2bb2o_1 _07693_ (.A1_N(_00892_),
    .A2_N(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .B2(_00979_),
    .X(_03078_));
 sky130_fd_sc_hd__nand2_1 _07694_ (.A(_00892_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ),
    .Y(_03079_));
 sky130_fd_sc_hd__a21bo_1 _07695_ (.A1(_03078_),
    .A2(_03079_),
    .B1_N(_03077_),
    .X(_03080_));
 sky130_fd_sc_hd__nand3_1 _07696_ (.A(_00891_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ),
    .C(_03075_),
    .Y(_03081_));
 sky130_fd_sc_hd__a31o_1 _07697_ (.A1(_03074_),
    .A2(_03080_),
    .A3(_03081_),
    .B1(_03073_),
    .X(_03082_));
 sky130_fd_sc_hd__and2b_1 _07698_ (.A_N(_03072_),
    .B(_03082_),
    .X(_03083_));
 sky130_fd_sc_hd__nand2_1 _07699_ (.A(_00886_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ),
    .Y(_03084_));
 sky130_fd_sc_hd__nor2_1 _07700_ (.A(_00888_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ),
    .Y(_03085_));
 sky130_fd_sc_hd__nor2_1 _07701_ (.A(_00886_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ),
    .Y(_03086_));
 sky130_fd_sc_hd__o21ai_1 _07702_ (.A1(_00887_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ),
    .B1(_03084_),
    .Y(_03087_));
 sky130_fd_sc_hd__a211o_1 _07703_ (.A1(_00887_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ),
    .B1(_03086_),
    .C1(_03087_),
    .X(_03088_));
 sky130_fd_sc_hd__or3_1 _07704_ (.A(_03083_),
    .B(_03085_),
    .C(_03088_),
    .X(_03089_));
 sky130_fd_sc_hd__or3b_1 _07705_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ),
    .B(_03086_),
    .C_N(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ),
    .X(_03090_));
 sky130_fd_sc_hd__a31o_1 _07706_ (.A1(_03084_),
    .A2(_03089_),
    .A3(_03090_),
    .B1(_03071_),
    .X(_03091_));
 sky130_fd_sc_hd__a32o_1 _07707_ (.A1(_03062_),
    .A2(_03064_),
    .A3(_03066_),
    .B1(_03061_),
    .B2(_03060_),
    .X(_03092_));
 sky130_fd_sc_hd__a21oi_1 _07708_ (.A1(_03068_),
    .A2(_03092_),
    .B1(_03067_),
    .Y(_03093_));
 sky130_fd_sc_hd__o21ai_1 _07709_ (.A1(net727),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp0[15] ),
    .B1(_03055_),
    .Y(_03094_));
 sky130_fd_sc_hd__o211a_1 _07710_ (.A1(_03057_),
    .A2(_03093_),
    .B1(_03094_),
    .C1(_03091_),
    .X(_03095_));
 sky130_fd_sc_hd__or4b_1 _07711_ (.A(_03072_),
    .B(_03073_),
    .C(_03085_),
    .D_N(_03077_),
    .X(_03096_));
 sky130_fd_sc_hd__o21ai_1 _07712_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .A2(_00979_),
    .B1(_03079_),
    .Y(_03097_));
 sky130_fd_sc_hd__or4_1 _07713_ (.A(_03078_),
    .B(_03088_),
    .C(_03096_),
    .D(_03097_),
    .X(_03098_));
 sky130_fd_sc_hd__nor2_1 _07714_ (.A(_03071_),
    .B(_03098_),
    .Y(_03099_));
 sky130_fd_sc_hd__o32ai_4 _07715_ (.A1(\u_pwm.u_pwm_1.cfg_comp0_center ),
    .A2(_03095_),
    .A3(_03099_),
    .B1(_03052_),
    .B2(_03054_),
    .Y(_03100_));
 sky130_fd_sc_hd__or2_1 _07716_ (.A(net727),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[15] ),
    .X(_03101_));
 sky130_fd_sc_hd__a22o_1 _07717_ (.A1(net727),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[15] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[14] ),
    .B2(_00879_),
    .X(_03102_));
 sky130_fd_sc_hd__a22o_1 _07718_ (.A1(_00880_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[13] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[12] ),
    .B2(_00881_),
    .X(_03103_));
 sky130_fd_sc_hd__or2_1 _07719_ (.A(_00881_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[12] ),
    .X(_03104_));
 sky130_fd_sc_hd__a22o_1 _07720_ (.A1(_00884_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[9] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[8] ),
    .B2(_00885_),
    .X(_03105_));
 sky130_fd_sc_hd__nand2b_1 _07721_ (.A_N(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[11] ),
    .Y(_03106_));
 sky130_fd_sc_hd__nand2b_1 _07722_ (.A_N(\u_pwm.u_pwm_1.cfg_pwm_comp1[11] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .Y(_03107_));
 sky130_fd_sc_hd__o211a_1 _07723_ (.A1(_00883_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[10] ),
    .B1(_03106_),
    .C1(_03107_),
    .X(_03108_));
 sky130_fd_sc_hd__o221a_1 _07724_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .A2(_00983_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[9] ),
    .B2(_00884_),
    .C1(_03108_),
    .X(_03109_));
 sky130_fd_sc_hd__o21ai_1 _07725_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .A2(_00983_),
    .B1(_03106_),
    .Y(_03110_));
 sky130_fd_sc_hd__a22o_1 _07726_ (.A1(_03105_),
    .A2(_03109_),
    .B1(_03110_),
    .B2(_03107_),
    .X(_03111_));
 sky130_fd_sc_hd__a21o_1 _07727_ (.A1(_03104_),
    .A2(_03111_),
    .B1(_03103_),
    .X(_03112_));
 sky130_fd_sc_hd__or2_1 _07728_ (.A(_00879_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[14] ),
    .X(_03113_));
 sky130_fd_sc_hd__or2_1 _07729_ (.A(_00880_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[13] ),
    .X(_03114_));
 sky130_fd_sc_hd__a31o_1 _07730_ (.A1(_03112_),
    .A2(_03113_),
    .A3(_03114_),
    .B1(_03102_),
    .X(_03115_));
 sky130_fd_sc_hd__a22o_1 _07731_ (.A1(_00886_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[6] ),
    .B2(_00887_),
    .X(_03116_));
 sky130_fd_sc_hd__or2_1 _07732_ (.A(net726),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[5] ),
    .X(_03117_));
 sky130_fd_sc_hd__a22o_1 _07733_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[4] ),
    .B2(_00889_),
    .X(_03118_));
 sky130_fd_sc_hd__nand2b_1 _07734_ (.A_N(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[1] ),
    .Y(_03119_));
 sky130_fd_sc_hd__nand2b_1 _07735_ (.A_N(\u_pwm.u_pwm_1.cfg_pwm_comp1[1] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .Y(_03120_));
 sky130_fd_sc_hd__o211ai_1 _07736_ (.A1(_00893_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[0] ),
    .B1(_03119_),
    .C1(_03120_),
    .Y(_03121_));
 sky130_fd_sc_hd__o2bb2a_1 _07737_ (.A1_N(_03119_),
    .A2_N(_03121_),
    .B1(_00891_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .X(_03122_));
 sky130_fd_sc_hd__a22o_1 _07738_ (.A1(_00890_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .B2(_00891_),
    .X(_03123_));
 sky130_fd_sc_hd__or2_1 _07739_ (.A(_00890_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ),
    .X(_03124_));
 sky130_fd_sc_hd__o21ba_1 _07740_ (.A1(_00889_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[4] ),
    .B1_N(_03118_),
    .X(_03125_));
 sky130_fd_sc_hd__o211a_1 _07741_ (.A1(_03122_),
    .A2(_03123_),
    .B1(_03125_),
    .C1(_03117_),
    .X(_03126_));
 sky130_fd_sc_hd__a22o_1 _07742_ (.A1(_03117_),
    .A2(_03118_),
    .B1(_03124_),
    .B2(_03126_),
    .X(_03127_));
 sky130_fd_sc_hd__or2_1 _07743_ (.A(_00887_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[6] ),
    .X(_03128_));
 sky130_fd_sc_hd__a21o_1 _07744_ (.A1(_03127_),
    .A2(_03128_),
    .B1(_03116_),
    .X(_03129_));
 sky130_fd_sc_hd__o211a_1 _07745_ (.A1(_00885_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp1[8] ),
    .B1(_03104_),
    .C1(_03114_),
    .X(_03130_));
 sky130_fd_sc_hd__and4bb_1 _07746_ (.A_N(_03103_),
    .B_N(_03105_),
    .C(_03113_),
    .D(_03130_),
    .X(_03131_));
 sky130_fd_sc_hd__and4b_1 _07747_ (.A_N(_03102_),
    .B(_03109_),
    .C(_03131_),
    .D(_03101_),
    .X(_03132_));
 sky130_fd_sc_hd__or2_1 _07748_ (.A(_00886_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ),
    .X(_03133_));
 sky130_fd_sc_hd__a32o_1 _07749_ (.A1(_03129_),
    .A2(_03132_),
    .A3(_03133_),
    .B1(_03115_),
    .B2(_03101_),
    .X(_03134_));
 sky130_fd_sc_hd__or4bb_1 _07750_ (.A(_03116_),
    .B(_03123_),
    .C_N(_03124_),
    .D_N(_03128_),
    .X(_03135_));
 sky130_fd_sc_hd__o221ai_1 _07751_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .A2(_00982_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .B2(_00891_),
    .C1(_03133_),
    .Y(_03136_));
 sky130_fd_sc_hd__nor2_1 _07752_ (.A(_03121_),
    .B(_03136_),
    .Y(_03137_));
 sky130_fd_sc_hd__and4b_1 _07753_ (.A_N(_03135_),
    .B(_03117_),
    .C(_03125_),
    .D(_03137_),
    .X(_03138_));
 sky130_fd_sc_hd__a21boi_1 _07754_ (.A1(_03132_),
    .A2(_03138_),
    .B1_N(_03134_),
    .Y(_03139_));
 sky130_fd_sc_hd__a22o_1 _07755_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[13] ),
    .A2(_03007_),
    .B1(_03008_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[12] ),
    .X(_03140_));
 sky130_fd_sc_hd__or2_1 _07756_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[11] ),
    .B(_03015_),
    .X(_03141_));
 sky130_fd_sc_hd__a22o_1 _07757_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[10] ),
    .A2(_03011_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[11] ),
    .X(_03142_));
 sky130_fd_sc_hd__a22o_1 _07758_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[8] ),
    .A2(_03006_),
    .B1(_03010_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[9] ),
    .X(_03143_));
 sky130_fd_sc_hd__o22a_1 _07759_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[9] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[10] ),
    .X(_03144_));
 sky130_fd_sc_hd__a21o_1 _07760_ (.A1(_03143_),
    .A2(_03144_),
    .B1(_03142_),
    .X(_03145_));
 sky130_fd_sc_hd__a22oi_1 _07761_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[6] ),
    .A2(_03026_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ),
    .Y(_03146_));
 sky130_fd_sc_hd__a22o_1 _07762_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[4] ),
    .A2(_03030_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[5] ),
    .X(_03147_));
 sky130_fd_sc_hd__a22o_1 _07763_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .A2(net588),
    .B1(net587),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ),
    .X(_03148_));
 sky130_fd_sc_hd__and2_1 _07764_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[1] ),
    .B(_03022_),
    .X(_03149_));
 sky130_fd_sc_hd__o22a_1 _07765_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[0] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[1] ),
    .X(_03150_));
 sky130_fd_sc_hd__o22a_1 _07766_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .A2(net588),
    .B1(_03149_),
    .B2(_03150_),
    .X(_03151_));
 sky130_fd_sc_hd__or2_1 _07767_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[4] ),
    .B(_03030_),
    .X(_03152_));
 sky130_fd_sc_hd__o21a_1 _07768_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[8] ),
    .A2(_03006_),
    .B1(_03141_),
    .X(_03153_));
 sky130_fd_sc_hd__and4bb_1 _07769_ (.A_N(_03142_),
    .B_N(_03143_),
    .C(_03144_),
    .D(_03153_),
    .X(_03154_));
 sky130_fd_sc_hd__o22a_1 _07770_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[6] ),
    .A2(_03026_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ),
    .X(_03155_));
 sky130_fd_sc_hd__o211a_1 _07771_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[5] ),
    .A2(_03031_),
    .B1(_03146_),
    .C1(_03155_),
    .X(_03156_));
 sky130_fd_sc_hd__and3b_1 _07772_ (.A_N(_03147_),
    .B(_03152_),
    .C(_03156_),
    .X(_03157_));
 sky130_fd_sc_hd__o22a_1 _07773_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ),
    .A2(net587),
    .B1(_03148_),
    .B2(_03151_),
    .X(_03158_));
 sky130_fd_sc_hd__o21ba_1 _07774_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ),
    .A2(_03027_),
    .B1_N(_03146_),
    .X(_03159_));
 sky130_fd_sc_hd__a221o_1 _07775_ (.A1(_03147_),
    .A2(_03156_),
    .B1(_03157_),
    .B2(_03158_),
    .C1(_03159_),
    .X(_03160_));
 sky130_fd_sc_hd__a22o_1 _07776_ (.A1(_03141_),
    .A2(_03145_),
    .B1(_03154_),
    .B2(_03160_),
    .X(_03161_));
 sky130_fd_sc_hd__or2_1 _07777_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[12] ),
    .B(_03008_),
    .X(_03162_));
 sky130_fd_sc_hd__nand2_1 _07778_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp1[0] ),
    .B(_03021_),
    .Y(_03163_));
 sky130_fd_sc_hd__o21ba_1 _07779_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ),
    .A2(net587),
    .B1_N(_03148_),
    .X(_03164_));
 sky130_fd_sc_hd__and4b_1 _07780_ (.A_N(_03149_),
    .B(_03150_),
    .C(_03154_),
    .D(_03164_),
    .X(_03165_));
 sky130_fd_sc_hd__o2111ai_2 _07781_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ),
    .A2(net588),
    .B1(_03157_),
    .C1(_03163_),
    .D1(_03165_),
    .Y(_03166_));
 sky130_fd_sc_hd__a31o_1 _07782_ (.A1(_03161_),
    .A2(_03162_),
    .A3(_03166_),
    .B1(_03140_),
    .X(_03167_));
 sky130_fd_sc_hd__o221a_1 _07783_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[14] ),
    .A2(_03004_),
    .B1(_03007_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp1[13] ),
    .C1(_03167_),
    .X(_03168_));
 sky130_fd_sc_hd__a211o_1 _07784_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp1[14] ),
    .A2(_03004_),
    .B1(_00984_),
    .C1(\u_pwm.u_pwm_1.cfg_pwm_comp1[15] ),
    .X(_03169_));
 sky130_fd_sc_hd__o22a_1 _07785_ (.A1(\u_pwm.u_pwm_1.cfg_comp1_center ),
    .A2(_03139_),
    .B1(_03168_),
    .B2(_03169_),
    .X(_03170_));
 sky130_fd_sc_hd__xnor2_1 _07786_ (.A(_03100_),
    .B(_03170_),
    .Y(_03171_));
 sky130_fd_sc_hd__a22o_1 _07787_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ),
    .A2(_03007_),
    .B1(_03008_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ),
    .X(_03172_));
 sky130_fd_sc_hd__a22o_1 _07788_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[8] ),
    .A2(_03006_),
    .B1(_03010_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ),
    .X(_03173_));
 sky130_fd_sc_hd__a22o_1 _07789_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[10] ),
    .A2(_03011_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[11] ),
    .X(_03174_));
 sky130_fd_sc_hd__o22a_1 _07790_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[10] ),
    .X(_03175_));
 sky130_fd_sc_hd__or4b_1 _07791_ (.A(_03172_),
    .B(_03173_),
    .C(_03174_),
    .D_N(_03175_),
    .X(_03176_));
 sky130_fd_sc_hd__o22a_1 _07792_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[14] ),
    .A2(_03004_),
    .B1(_03007_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ),
    .X(_03177_));
 sky130_fd_sc_hd__o221ai_1 _07793_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ),
    .A2(_03008_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[11] ),
    .C1(_03177_),
    .Y(_03178_));
 sky130_fd_sc_hd__a21o_1 _07794_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[14] ),
    .A2(_03004_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[15] ),
    .X(_03179_));
 sky130_fd_sc_hd__o22a_1 _07795_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[8] ),
    .A2(_03006_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ),
    .X(_03180_));
 sky130_fd_sc_hd__or4b_1 _07796_ (.A(_03176_),
    .B(_03178_),
    .C(_03179_),
    .D_N(_03180_),
    .X(_03181_));
 sky130_fd_sc_hd__a22o_1 _07797_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ),
    .A2(_03026_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ),
    .X(_03182_));
 sky130_fd_sc_hd__o22a_1 _07798_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ),
    .A2(_03026_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ),
    .X(_03183_));
 sky130_fd_sc_hd__a22o_1 _07799_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ),
    .A2(_03030_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ),
    .X(_03184_));
 sky130_fd_sc_hd__o22a_1 _07800_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ),
    .A2(_03030_),
    .B1(net587),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ),
    .X(_03185_));
 sky130_fd_sc_hd__a22o_1 _07801_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ),
    .A2(net588),
    .B1(net587),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ),
    .X(_03186_));
 sky130_fd_sc_hd__nor2_1 _07802_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ),
    .B(net588),
    .Y(_03187_));
 sky130_fd_sc_hd__nand2_1 _07803_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ),
    .B(_03022_),
    .Y(_03188_));
 sky130_fd_sc_hd__o22a_1 _07804_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ),
    .X(_03189_));
 sky130_fd_sc_hd__nand2_1 _07805_ (.A(_03188_),
    .B(_03189_),
    .Y(_03190_));
 sky130_fd_sc_hd__a21oi_1 _07806_ (.A1(_03188_),
    .A2(_03190_),
    .B1(_03187_),
    .Y(_03191_));
 sky130_fd_sc_hd__o21a_1 _07807_ (.A1(_03186_),
    .A2(_03191_),
    .B1(_03185_),
    .X(_03192_));
 sky130_fd_sc_hd__o21a_1 _07808_ (.A1(_03184_),
    .A2(_03192_),
    .B1(_03183_),
    .X(_03193_));
 sky130_fd_sc_hd__o21ba_1 _07809_ (.A1(_03182_),
    .A2(_03193_),
    .B1_N(_03181_),
    .X(_03194_));
 sky130_fd_sc_hd__a21oi_1 _07810_ (.A1(_03173_),
    .A2(_03175_),
    .B1(_03174_),
    .Y(_03195_));
 sky130_fd_sc_hd__nor2_1 _07811_ (.A(_03178_),
    .B(_03195_),
    .Y(_03196_));
 sky130_fd_sc_hd__a2111o_1 _07812_ (.A1(_03172_),
    .A2(_03177_),
    .B1(_03179_),
    .C1(_03194_),
    .D1(_03196_),
    .X(_03197_));
 sky130_fd_sc_hd__nand2_1 _07813_ (.A(_03183_),
    .B(_03185_),
    .Y(_03198_));
 sky130_fd_sc_hd__or3_1 _07814_ (.A(_03184_),
    .B(_03186_),
    .C(_03198_),
    .X(_03199_));
 sky130_fd_sc_hd__a211o_1 _07815_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ),
    .A2(_03021_),
    .B1(_03182_),
    .C1(_03187_),
    .X(_03200_));
 sky130_fd_sc_hd__or4_1 _07816_ (.A(_03181_),
    .B(_03190_),
    .C(_03199_),
    .D(_03200_),
    .X(_03201_));
 sky130_fd_sc_hd__nor2_1 _07817_ (.A(_00878_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp2[15] ),
    .Y(_03202_));
 sky130_fd_sc_hd__o22a_1 _07818_ (.A1(_00884_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[10] ),
    .B2(_00883_),
    .X(_03203_));
 sky130_fd_sc_hd__a22o_1 _07819_ (.A1(_00885_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[8] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ),
    .B2(_00884_),
    .X(_03204_));
 sky130_fd_sc_hd__nand2_1 _07820_ (.A(_03203_),
    .B(_03204_),
    .Y(_03205_));
 sky130_fd_sc_hd__o221a_1 _07821_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .A2(_00962_),
    .B1(_00963_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .C1(_03205_),
    .X(_03206_));
 sky130_fd_sc_hd__a2bb2o_1 _07822_ (.A1_N(_00881_),
    .A2_N(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .B2(_00963_),
    .X(_03207_));
 sky130_fd_sc_hd__a22o_1 _07823_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .A2(_00964_),
    .B1(_00965_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .X(_03208_));
 sky130_fd_sc_hd__a22o_1 _07824_ (.A1(_00879_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[14] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[15] ),
    .B2(net727),
    .X(_03209_));
 sky130_fd_sc_hd__a22o_1 _07825_ (.A1(_00881_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ),
    .B2(_00880_),
    .X(_03210_));
 sky130_fd_sc_hd__o21ba_1 _07826_ (.A1(_03206_),
    .A2(_03207_),
    .B1_N(_03210_),
    .X(_03211_));
 sky130_fd_sc_hd__a221o_1 _07827_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .A2(_00964_),
    .B1(_00965_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .C1(_03211_),
    .X(_03212_));
 sky130_fd_sc_hd__and2b_1 _07828_ (.A_N(_03209_),
    .B(_03212_),
    .X(_03213_));
 sky130_fd_sc_hd__a22o_1 _07829_ (.A1(_00887_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ),
    .B2(_00886_),
    .X(_03214_));
 sky130_fd_sc_hd__a22o_1 _07830_ (.A1(_00889_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ),
    .B2(net726),
    .X(_03215_));
 sky130_fd_sc_hd__o22a_1 _07831_ (.A1(_00890_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ),
    .B2(_00889_),
    .X(_03216_));
 sky130_fd_sc_hd__nor2_1 _07832_ (.A(_00891_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ),
    .Y(_03217_));
 sky130_fd_sc_hd__nand2_1 _07833_ (.A(_00892_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ),
    .Y(_03218_));
 sky130_fd_sc_hd__o22a_1 _07834_ (.A1(_00893_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ),
    .B2(_00892_),
    .X(_03219_));
 sky130_fd_sc_hd__nand2_1 _07835_ (.A(_03218_),
    .B(_03219_),
    .Y(_03220_));
 sky130_fd_sc_hd__a21oi_1 _07836_ (.A1(_03218_),
    .A2(_03220_),
    .B1(_03217_),
    .Y(_03221_));
 sky130_fd_sc_hd__a22o_1 _07837_ (.A1(_00891_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ),
    .B2(_00890_),
    .X(_03222_));
 sky130_fd_sc_hd__o21a_1 _07838_ (.A1(_03221_),
    .A2(_03222_),
    .B1(_03216_),
    .X(_03223_));
 sky130_fd_sc_hd__o22ai_1 _07839_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ),
    .B2(_00887_),
    .Y(_03224_));
 sky130_fd_sc_hd__o21ba_1 _07840_ (.A1(_03215_),
    .A2(_03223_),
    .B1_N(_03224_),
    .X(_03225_));
 sky130_fd_sc_hd__nor2_1 _07841_ (.A(_03214_),
    .B(_03225_),
    .Y(_03226_));
 sky130_fd_sc_hd__o221a_1 _07842_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .A2(_00962_),
    .B1(_00963_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .C1(_03203_),
    .X(_03227_));
 sky130_fd_sc_hd__nor2_1 _07843_ (.A(_00886_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ),
    .Y(_03228_));
 sky130_fd_sc_hd__or3b_1 _07844_ (.A(_03204_),
    .B(_03210_),
    .C_N(_03227_),
    .X(_03229_));
 sky130_fd_sc_hd__a211o_1 _07845_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ),
    .A2(_00961_),
    .B1(_03207_),
    .C1(_03208_),
    .X(_03230_));
 sky130_fd_sc_hd__or4_1 _07846_ (.A(_03202_),
    .B(_03209_),
    .C(_03229_),
    .D(_03230_),
    .X(_03231_));
 sky130_fd_sc_hd__o32a_1 _07847_ (.A1(_03226_),
    .A2(_03228_),
    .A3(_03231_),
    .B1(_03213_),
    .B2(_03202_),
    .X(_03232_));
 sky130_fd_sc_hd__a221o_1 _07848_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .A2(_00959_),
    .B1(_00960_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .C1(_03222_),
    .X(_03233_));
 sky130_fd_sc_hd__a2111o_1 _07849_ (.A1(_00893_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ),
    .B1(_03214_),
    .C1(_03217_),
    .D1(_03220_),
    .X(_03234_));
 sky130_fd_sc_hd__or4_1 _07850_ (.A(_03215_),
    .B(_03224_),
    .C(_03233_),
    .D(_03234_),
    .X(_03235_));
 sky130_fd_sc_hd__nor3_1 _07851_ (.A(_03228_),
    .B(_03231_),
    .C(_03235_),
    .Y(_03236_));
 sky130_fd_sc_hd__nor3_1 _07852_ (.A(\u_pwm.u_pwm_1.cfg_comp2_center ),
    .B(_03232_),
    .C(_03236_),
    .Y(_03237_));
 sky130_fd_sc_hd__a31o_1 _07853_ (.A1(\u_pwm.u_pwm_1.cfg_comp2_center ),
    .A2(_03197_),
    .A3(_03201_),
    .B1(_03237_),
    .X(_03238_));
 sky130_fd_sc_hd__xnor2_1 _07854_ (.A(_03171_),
    .B(_03238_),
    .Y(_03239_));
 sky130_fd_sc_hd__a22o_1 _07855_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ),
    .A2(_03026_),
    .B1(_03027_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ),
    .X(_03240_));
 sky130_fd_sc_hd__a22o_1 _07856_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .A2(_03030_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ),
    .X(_03241_));
 sky130_fd_sc_hd__a22o_1 _07857_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .A2(net588),
    .B1(net587),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .X(_03242_));
 sky130_fd_sc_hd__nand2_1 _07858_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .B(_03022_),
    .Y(_03243_));
 sky130_fd_sc_hd__o22a_1 _07859_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ),
    .A2(_03021_),
    .B1(_03022_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .X(_03244_));
 sky130_fd_sc_hd__nand2_1 _07860_ (.A(_03243_),
    .B(_03244_),
    .Y(_03245_));
 sky130_fd_sc_hd__o2bb2a_1 _07861_ (.A1_N(_03243_),
    .A2_N(_03245_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .B2(net588),
    .X(_03246_));
 sky130_fd_sc_hd__nor2_1 _07862_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .B(_03030_),
    .Y(_03247_));
 sky130_fd_sc_hd__or2_1 _07863_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .B(net587),
    .X(_03248_));
 sky130_fd_sc_hd__o221a_1 _07864_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .A2(_03030_),
    .B1(_03242_),
    .B2(_03246_),
    .C1(_03248_),
    .X(_03249_));
 sky130_fd_sc_hd__o22a_1 _07865_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ),
    .A2(_03026_),
    .B1(_03031_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ),
    .X(_03250_));
 sky130_fd_sc_hd__o21a_1 _07866_ (.A1(_03241_),
    .A2(_03249_),
    .B1(_03250_),
    .X(_03251_));
 sky130_fd_sc_hd__nor2_1 _07867_ (.A(_03240_),
    .B(_03251_),
    .Y(_03252_));
 sky130_fd_sc_hd__a22o_1 _07868_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .A2(_03011_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[11] ),
    .X(_03253_));
 sky130_fd_sc_hd__a22o_1 _07869_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[13] ),
    .A2(_03007_),
    .B1(_03008_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[12] ),
    .X(_03254_));
 sky130_fd_sc_hd__o22a_1 _07870_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[12] ),
    .A2(_03008_),
    .B1(_03015_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[11] ),
    .X(_03255_));
 sky130_fd_sc_hd__a21o_1 _07871_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[14] ),
    .A2(_03004_),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ),
    .X(_03256_));
 sky130_fd_sc_hd__o22a_1 _07872_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[14] ),
    .A2(_03004_),
    .B1(_03007_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[13] ),
    .X(_03257_));
 sky130_fd_sc_hd__a22o_1 _07873_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ),
    .A2(_03006_),
    .B1(_03010_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .X(_03258_));
 sky130_fd_sc_hd__o21ai_1 _07874_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ),
    .A2(_03006_),
    .B1(_03257_),
    .Y(_03259_));
 sky130_fd_sc_hd__o221a_1 _07875_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .C1(_03255_),
    .X(_03260_));
 sky130_fd_sc_hd__or3b_1 _07876_ (.A(_03253_),
    .B(_03258_),
    .C_N(_03260_),
    .X(_03261_));
 sky130_fd_sc_hd__or4_1 _07877_ (.A(_03254_),
    .B(_03256_),
    .C(_03259_),
    .D(_03261_),
    .X(_03262_));
 sky130_fd_sc_hd__nor2_1 _07878_ (.A(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ),
    .B(_03027_),
    .Y(_03263_));
 sky130_fd_sc_hd__or3_1 _07879_ (.A(_03252_),
    .B(_03262_),
    .C(_03263_),
    .X(_03264_));
 sky130_fd_sc_hd__o221a_1 _07880_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .A2(_03010_),
    .B1(_03011_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .C1(_03258_),
    .X(_03265_));
 sky130_fd_sc_hd__o21a_1 _07881_ (.A1(_03253_),
    .A2(_03265_),
    .B1(_03255_),
    .X(_03266_));
 sky130_fd_sc_hd__o21ai_1 _07882_ (.A1(_03254_),
    .A2(_03266_),
    .B1(_03257_),
    .Y(_03267_));
 sky130_fd_sc_hd__and3b_1 _07883_ (.A_N(_03256_),
    .B(_03264_),
    .C(_03267_),
    .X(_03268_));
 sky130_fd_sc_hd__o221ai_1 _07884_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .A2(_03038_),
    .B1(_03041_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .C1(_03250_),
    .Y(_03269_));
 sky130_fd_sc_hd__a2111o_1 _07885_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ),
    .A2(_03021_),
    .B1(_03247_),
    .C1(_03263_),
    .D1(_03269_),
    .X(_03270_));
 sky130_fd_sc_hd__or4_1 _07886_ (.A(_03240_),
    .B(_03241_),
    .C(_03242_),
    .D(_03262_),
    .X(_03271_));
 sky130_fd_sc_hd__o31ai_1 _07887_ (.A1(_03245_),
    .A2(_03270_),
    .A3(_03271_),
    .B1(\u_pwm.u_pwm_1.cfg_comp3_center ),
    .Y(_03272_));
 sky130_fd_sc_hd__nor2_1 _07888_ (.A(net727),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ),
    .Y(_03273_));
 sky130_fd_sc_hd__a22o_1 _07889_ (.A1(_00883_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[11] ),
    .B2(_00882_),
    .X(_03274_));
 sky130_fd_sc_hd__a22o_1 _07890_ (.A1(_00885_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .B2(_00884_),
    .X(_03275_));
 sky130_fd_sc_hd__o22a_1 _07891_ (.A1(_00884_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ),
    .B2(_00883_),
    .X(_03276_));
 sky130_fd_sc_hd__a21oi_1 _07892_ (.A1(_03275_),
    .A2(_03276_),
    .B1(_03274_),
    .Y(_03277_));
 sky130_fd_sc_hd__a22o_1 _07893_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .A2(_00969_),
    .B1(_00970_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .X(_03278_));
 sky130_fd_sc_hd__a221o_1 _07894_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ),
    .A2(_00967_),
    .B1(_00968_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .C1(_03278_),
    .X(_03279_));
 sky130_fd_sc_hd__o2bb2a_1 _07895_ (.A1_N(net727),
    .A2_N(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ),
    .B2(_00970_),
    .X(_03280_));
 sky130_fd_sc_hd__o22a_1 _07896_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .A2(_00968_),
    .B1(_00969_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .X(_03281_));
 sky130_fd_sc_hd__o221a_1 _07897_ (.A1(_03277_),
    .A2(_03279_),
    .B1(_03281_),
    .B2(_03278_),
    .C1(_03280_),
    .X(_03282_));
 sky130_fd_sc_hd__a22o_1 _07898_ (.A1(_00887_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ),
    .B2(_00886_),
    .X(_03283_));
 sky130_fd_sc_hd__a22o_1 _07899_ (.A1(_00889_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ),
    .B2(net726),
    .X(_03284_));
 sky130_fd_sc_hd__o22ai_1 _07900_ (.A1(_00890_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ),
    .B2(_00889_),
    .Y(_03285_));
 sky130_fd_sc_hd__nand2_1 _07901_ (.A(_00892_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .Y(_03286_));
 sky130_fd_sc_hd__o22ai_1 _07902_ (.A1(_00893_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .B2(_00892_),
    .Y(_03287_));
 sky130_fd_sc_hd__o2bb2a_1 _07903_ (.A1_N(_03286_),
    .A2_N(_03287_),
    .B1(_00891_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .X(_03288_));
 sky130_fd_sc_hd__a22o_1 _07904_ (.A1(_00891_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ),
    .B2(_00890_),
    .X(_03289_));
 sky130_fd_sc_hd__o21ba_1 _07905_ (.A1(_03288_),
    .A2(_03289_),
    .B1_N(_03285_),
    .X(_03290_));
 sky130_fd_sc_hd__o22a_1 _07906_ (.A1(net726),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ),
    .B2(_00887_),
    .X(_03291_));
 sky130_fd_sc_hd__o21a_1 _07907_ (.A1(_03284_),
    .A2(_03290_),
    .B1(_03291_),
    .X(_03292_));
 sky130_fd_sc_hd__nor2_1 _07908_ (.A(_03283_),
    .B(_03292_),
    .Y(_03293_));
 sky130_fd_sc_hd__nor2_1 _07909_ (.A(_00886_),
    .B(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ),
    .Y(_03294_));
 sky130_fd_sc_hd__o221a_1 _07910_ (.A1(_00885_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ),
    .B2(net727),
    .C1(_03280_),
    .X(_03295_));
 sky130_fd_sc_hd__and4bb_1 _07911_ (.A_N(_03274_),
    .B_N(_03275_),
    .C(_03276_),
    .D(_03281_),
    .X(_03296_));
 sky130_fd_sc_hd__or4bb_1 _07912_ (.A(_03279_),
    .B(_03294_),
    .C_N(_03295_),
    .D_N(_03296_),
    .X(_03297_));
 sky130_fd_sc_hd__o22a_1 _07913_ (.A1(_03273_),
    .A2(_03282_),
    .B1(_03293_),
    .B2(_03297_),
    .X(_03298_));
 sky130_fd_sc_hd__or4b_1 _07914_ (.A(_03284_),
    .B(_03285_),
    .C(_03287_),
    .D_N(_03291_),
    .X(_03299_));
 sky130_fd_sc_hd__a221o_1 _07915_ (.A1(_00892_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ),
    .B1(_00966_),
    .B2(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ),
    .C1(_03283_),
    .X(_03300_));
 sky130_fd_sc_hd__a2111o_1 _07916_ (.A1(_00893_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ),
    .B1(_03289_),
    .C1(_03299_),
    .D1(_03300_),
    .X(_03301_));
 sky130_fd_sc_hd__nor2_1 _07917_ (.A(_03297_),
    .B(_03301_),
    .Y(_03302_));
 sky130_fd_sc_hd__o32a_1 _07918_ (.A1(\u_pwm.u_pwm_1.cfg_comp3_center ),
    .A2(_03298_),
    .A3(_03302_),
    .B1(_03268_),
    .B2(_03272_),
    .X(_03303_));
 sky130_fd_sc_hd__xnor2_1 _07919_ (.A(_03239_),
    .B(_03303_),
    .Y(_03304_));
 sky130_fd_sc_hd__nor2_1 _07920_ (.A(\u_pwm.u_pwm_1.cfg_pwm_mode[1] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_mode[0] ),
    .Y(_03305_));
 sky130_fd_sc_hd__or3_1 _07921_ (.A(\u_pwm.u_pwm_1.cfg_pwm_mode[1] ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_mode[0] ),
    .C(_03100_),
    .X(_03306_));
 sky130_fd_sc_hd__o22a_1 _07922_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_mode[1] ),
    .A2(_03171_),
    .B1(_03239_),
    .B2(\u_pwm.u_pwm_1.cfg_pwm_mode[0] ),
    .X(_03307_));
 sky130_fd_sc_hd__o21ai_1 _07923_ (.A1(_03305_),
    .A2(_03307_),
    .B1(_03306_),
    .Y(_03308_));
 sky130_fd_sc_hd__a31o_1 _07924_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_mode[1] ),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_mode[0] ),
    .A3(_03304_),
    .B1(_03308_),
    .X(\u_pwm.u_pwm_1.u_pwm.pwm_wfm_i ));
 sky130_fd_sc_hd__and3_1 _07925_ (.A(net1355),
    .B(net1372),
    .C(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ),
    .X(_03309_));
 sky130_fd_sc_hd__a221o_1 _07926_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .A2(net1244),
    .B1(net1158),
    .B2(net1824),
    .C1(_03309_),
    .X(\u_pwm.u_glbl_reg.reg_out[0] ));
 sky130_fd_sc_hd__and3_1 _07927_ (.A(net1355),
    .B(net1372),
    .C(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ),
    .X(_03310_));
 sky130_fd_sc_hd__a221o_1 _07928_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .A2(net1244),
    .B1(net1158),
    .B2(net1822),
    .C1(_03310_),
    .X(\u_pwm.u_glbl_reg.reg_out[1] ));
 sky130_fd_sc_hd__and3_1 _07929_ (.A(net1355),
    .B(net1372),
    .C(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(_03311_));
 sky130_fd_sc_hd__a221o_1 _07930_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .A2(net1239),
    .B1(net1157),
    .B2(net1834),
    .C1(_03311_),
    .X(\u_pwm.u_glbl_reg.reg_out[2] ));
 sky130_fd_sc_hd__and3_1 _07931_ (.A(net1354),
    .B(net1261),
    .C(net1976),
    .X(\u_pwm.u_glbl_reg.reg_out[3] ));
 sky130_fd_sc_hd__and3_1 _07932_ (.A(net1354),
    .B(net1261),
    .C(net1977),
    .X(\u_pwm.u_glbl_reg.reg_out[4] ));
 sky130_fd_sc_hd__and3_1 _07933_ (.A(net1356),
    .B(net1261),
    .C(net1970),
    .X(\u_pwm.u_glbl_reg.reg_out[5] ));
 sky130_fd_sc_hd__and2_1 _07934_ (.A(net1948),
    .B(net1243),
    .X(\u_pwm.u_glbl_reg.reg_out[8] ));
 sky130_fd_sc_hd__and2_1 _07935_ (.A(net1816),
    .B(net1239),
    .X(\u_pwm.u_glbl_reg.reg_out[9] ));
 sky130_fd_sc_hd__and2_1 _07936_ (.A(net1826),
    .B(net1239),
    .X(\u_pwm.u_glbl_reg.reg_out[10] ));
 sky130_fd_sc_hd__and2_1 _07937_ (.A(net2016),
    .B(net1243),
    .X(\u_pwm.u_glbl_reg.reg_out[16] ));
 sky130_fd_sc_hd__and2_1 _07938_ (.A(net2007),
    .B(net1239),
    .X(\u_pwm.u_glbl_reg.reg_out[17] ));
 sky130_fd_sc_hd__and2_1 _07939_ (.A(net2046),
    .B(net1243),
    .X(\u_pwm.u_glbl_reg.reg_out[18] ));
 sky130_fd_sc_hd__a221o_1 _07940_ (.A1(net1264),
    .A2(\u_timer.cfg_timer1[0] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[0] ),
    .C1(net1250),
    .X(_03312_));
 sky130_fd_sc_hd__and3_1 _07941_ (.A(net1283),
    .B(net1370),
    .C(\u_timer.cfg_timer0[0] ),
    .X(_03313_));
 sky130_fd_sc_hd__o22a_1 _07942_ (.A1(\u_timer.cfg_pulse_1us[0] ),
    .A2(net1231),
    .B1(_03312_),
    .B2(_03313_),
    .X(\u_timer.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__and3_1 _07943_ (.A(net1283),
    .B(net1370),
    .C(\u_timer.cfg_timer0[1] ),
    .X(_03314_));
 sky130_fd_sc_hd__a221o_1 _07944_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[1] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[1] ),
    .C1(net1250),
    .X(_03315_));
 sky130_fd_sc_hd__o22a_1 _07945_ (.A1(\u_timer.cfg_pulse_1us[1] ),
    .A2(net1231),
    .B1(_03314_),
    .B2(_03315_),
    .X(\u_timer.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__a221o_1 _07946_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[2] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[2] ),
    .C1(net1250),
    .X(_03316_));
 sky130_fd_sc_hd__and3_1 _07947_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[2] ),
    .X(_03317_));
 sky130_fd_sc_hd__o22a_2 _07948_ (.A1(\u_timer.cfg_pulse_1us[2] ),
    .A2(net1231),
    .B1(_03316_),
    .B2(_03317_),
    .X(\u_timer.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__a221o_1 _07949_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[3] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[3] ),
    .C1(net1250),
    .X(_03318_));
 sky130_fd_sc_hd__and3_1 _07950_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[3] ),
    .X(_03319_));
 sky130_fd_sc_hd__o22a_2 _07951_ (.A1(\u_timer.cfg_pulse_1us[3] ),
    .A2(net1231),
    .B1(_03318_),
    .B2(_03319_),
    .X(\u_timer.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__a221o_1 _07952_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[4] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[4] ),
    .C1(net1251),
    .X(_03320_));
 sky130_fd_sc_hd__and3_1 _07953_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[4] ),
    .X(_03321_));
 sky130_fd_sc_hd__o22a_1 _07954_ (.A1(\u_timer.cfg_pulse_1us[4] ),
    .A2(net1231),
    .B1(_03320_),
    .B2(_03321_),
    .X(\u_timer.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__a221o_1 _07955_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[5] ),
    .B1(net1149),
    .B2(\u_timer.cfg_timer2[5] ),
    .C1(net1251),
    .X(_03322_));
 sky130_fd_sc_hd__and3_1 _07956_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[5] ),
    .X(_03323_));
 sky130_fd_sc_hd__o22a_1 _07957_ (.A1(\u_timer.cfg_pulse_1us[5] ),
    .A2(net1232),
    .B1(_03322_),
    .B2(_03323_),
    .X(\u_timer.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__and3_1 _07958_ (.A(net1283),
    .B(net1371),
    .C(\u_timer.cfg_timer0[6] ),
    .X(_03324_));
 sky130_fd_sc_hd__a221o_1 _07959_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[6] ),
    .B1(net1149),
    .B2(\u_timer.cfg_timer2[6] ),
    .C1(net1251),
    .X(_03325_));
 sky130_fd_sc_hd__o22a_1 _07960_ (.A1(\u_timer.cfg_pulse_1us[6] ),
    .A2(net1232),
    .B1(_03324_),
    .B2(_03325_),
    .X(\u_timer.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__and3_1 _07961_ (.A(net1282),
    .B(net1371),
    .C(\u_timer.cfg_timer0[7] ),
    .X(_03326_));
 sky130_fd_sc_hd__a221o_1 _07962_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[7] ),
    .B1(net1149),
    .B2(\u_timer.cfg_timer2[7] ),
    .C1(net1251),
    .X(_03327_));
 sky130_fd_sc_hd__o22a_1 _07963_ (.A1(\u_timer.cfg_pulse_1us[7] ),
    .A2(net1231),
    .B1(_03326_),
    .B2(_03327_),
    .X(\u_timer.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__a221o_1 _07964_ (.A1(net1263),
    .A2(net2022),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[8] ),
    .C1(net1250),
    .X(_03328_));
 sky130_fd_sc_hd__and3_1 _07965_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[8] ),
    .X(_03329_));
 sky130_fd_sc_hd__o22a_1 _07966_ (.A1(\u_timer.cfg_pulse_1us[8] ),
    .A2(net1231),
    .B1(_03328_),
    .B2(_03329_),
    .X(\u_timer.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__a221o_1 _07967_ (.A1(net1263),
    .A2(net2021),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[9] ),
    .C1(net1250),
    .X(_03330_));
 sky130_fd_sc_hd__and3_1 _07968_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[9] ),
    .X(_03331_));
 sky130_fd_sc_hd__o22a_1 _07969_ (.A1(\u_timer.cfg_pulse_1us[9] ),
    .A2(net1231),
    .B1(_03330_),
    .B2(_03331_),
    .X(\u_timer.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__a221o_1 _07970_ (.A1(net1263),
    .A2(\u_timer.cfg_timer1[10] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[10] ),
    .C1(net1250),
    .X(_03332_));
 sky130_fd_sc_hd__and3_1 _07971_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[10] ),
    .X(_03333_));
 sky130_fd_sc_hd__o22a_1 _07972_ (.A1(net2335),
    .A2(net1231),
    .B1(_03332_),
    .B2(_03333_),
    .X(\u_timer.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__a221o_1 _07973_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[11] ),
    .B1(net1148),
    .B2(\u_timer.cfg_timer2[11] ),
    .C1(net1250),
    .X(_03334_));
 sky130_fd_sc_hd__and3_1 _07974_ (.A(net1282),
    .B(net1370),
    .C(\u_timer.cfg_timer0[11] ),
    .X(_03335_));
 sky130_fd_sc_hd__o22a_1 _07975_ (.A1(net2292),
    .A2(net1231),
    .B1(_03334_),
    .B2(_03335_),
    .X(\u_timer.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__and3_1 _07976_ (.A(net1282),
    .B(net1369),
    .C(\u_timer.cfg_timer0[12] ),
    .X(_03336_));
 sky130_fd_sc_hd__a221o_1 _07977_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[12] ),
    .B1(net1150),
    .B2(\u_timer.cfg_timer2[12] ),
    .C1(net1248),
    .X(_03337_));
 sky130_fd_sc_hd__o22a_1 _07978_ (.A1(net2294),
    .A2(net1232),
    .B1(_03336_),
    .B2(_03337_),
    .X(\u_timer.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__and3_1 _07979_ (.A(net1280),
    .B(net1369),
    .C(\u_timer.cfg_timer0[13] ),
    .X(_03338_));
 sky130_fd_sc_hd__a221o_1 _07980_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[13] ),
    .B1(net1150),
    .B2(\u_timer.cfg_timer2[13] ),
    .C1(net1248),
    .X(_03339_));
 sky130_fd_sc_hd__o22a_1 _07981_ (.A1(net2314),
    .A2(net1232),
    .B1(_03338_),
    .B2(_03339_),
    .X(\u_timer.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__and3_1 _07982_ (.A(net1280),
    .B(net1369),
    .C(\u_timer.cfg_timer0[14] ),
    .X(_03340_));
 sky130_fd_sc_hd__a221o_1 _07983_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[14] ),
    .B1(net1150),
    .B2(\u_timer.cfg_timer2[14] ),
    .C1(net1248),
    .X(_03341_));
 sky130_fd_sc_hd__o22a_1 _07984_ (.A1(net2268),
    .A2(net1232),
    .B1(_03340_),
    .B2(_03341_),
    .X(\u_timer.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__a221o_1 _07985_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[15] ),
    .B1(net1150),
    .B2(\u_timer.cfg_timer2[15] ),
    .C1(net1248),
    .X(_03342_));
 sky130_fd_sc_hd__and3_1 _07986_ (.A(net1280),
    .B(net1371),
    .C(\u_timer.cfg_timer0[15] ),
    .X(_03343_));
 sky130_fd_sc_hd__o22a_1 _07987_ (.A1(net2267),
    .A2(net1232),
    .B1(_03342_),
    .B2(_03343_),
    .X(\u_timer.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__a22o_1 _07988_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[16] ),
    .B1(net1150),
    .B2(\u_timer.cfg_timer2[16] ),
    .X(_03344_));
 sky130_fd_sc_hd__a21oi_1 _07989_ (.A1(net1369),
    .A2(_00848_),
    .B1(net1357),
    .Y(_03345_));
 sky130_fd_sc_hd__o22a_1 _07990_ (.A1(net2274),
    .A2(net1232),
    .B1(_03344_),
    .B2(_03345_),
    .X(\u_timer.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__a221o_1 _07991_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[17] ),
    .B1(\u_timer.cfg_timer2[17] ),
    .B2(net1150),
    .C1(net1248),
    .X(_03346_));
 sky130_fd_sc_hd__and3_1 _07992_ (.A(net1280),
    .B(net1369),
    .C(\u_timer.cfg_timer0[17] ),
    .X(_03347_));
 sky130_fd_sc_hd__o22a_1 _07993_ (.A1(net2296),
    .A2(net1232),
    .B1(_03346_),
    .B2(_03347_),
    .X(\u_timer.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__and3_1 _07994_ (.A(net1280),
    .B(net1369),
    .C(\u_timer.cfg_timer0[18] ),
    .X(_03348_));
 sky130_fd_sc_hd__a221o_1 _07995_ (.A1(net1262),
    .A2(\u_timer.cfg_timer1[18] ),
    .B1(\u_timer.cfg_timer2[18] ),
    .B2(net1150),
    .C1(net1248),
    .X(_03349_));
 sky130_fd_sc_hd__o22a_1 _07996_ (.A1(net2327),
    .A2(net1232),
    .B1(_03348_),
    .B2(_03349_),
    .X(\u_timer.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__o21a_1 _07997_ (.A1(net1260),
    .A2(\u_timer.u_reg.reg_1[19] ),
    .B1(net1275),
    .X(_03350_));
 sky130_fd_sc_hd__a22o_1 _07998_ (.A1(net1260),
    .A2(\u_timer.u_reg.reg_2[19] ),
    .B1(net1146),
    .B2(\u_timer.u_reg.reg_3[19] ),
    .X(_03351_));
 sky130_fd_sc_hd__o22a_1 _07999_ (.A1(net2338),
    .A2(net1227),
    .B1(_03350_),
    .B2(_03351_),
    .X(\u_timer.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__o21a_1 _08000_ (.A1(net1275),
    .A2(\u_timer.u_reg.reg_2[20] ),
    .B1(net1260),
    .X(_03352_));
 sky130_fd_sc_hd__a221o_1 _08001_ (.A1(net1275),
    .A2(\u_timer.u_reg.reg_1[20] ),
    .B1(net1146),
    .B2(\u_timer.u_reg.reg_3[20] ),
    .C1(_03352_),
    .X(_03353_));
 sky130_fd_sc_hd__o21a_1 _08002_ (.A1(net2284),
    .A2(net1227),
    .B1(_03353_),
    .X(\u_timer.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__o21a_1 _08003_ (.A1(net1280),
    .A2(\u_timer.u_reg.reg_2[21] ),
    .B1(net1262),
    .X(_03354_));
 sky130_fd_sc_hd__a221o_1 _08004_ (.A1(net1280),
    .A2(\u_timer.u_reg.reg_1[21] ),
    .B1(net1150),
    .B2(\u_timer.u_reg.reg_3[21] ),
    .C1(_03354_),
    .X(_03355_));
 sky130_fd_sc_hd__o21a_1 _08005_ (.A1(net2231),
    .A2(net1232),
    .B1(_03355_),
    .X(\u_timer.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__o21a_1 _08006_ (.A1(net1260),
    .A2(\u_timer.u_reg.reg_1[22] ),
    .B1(net1275),
    .X(_03356_));
 sky130_fd_sc_hd__a22o_1 _08007_ (.A1(net1260),
    .A2(\u_timer.u_reg.reg_2[22] ),
    .B1(net1146),
    .B2(\u_timer.u_reg.reg_3[22] ),
    .X(_03357_));
 sky130_fd_sc_hd__o22a_1 _08008_ (.A1(net2301),
    .A2(net1227),
    .B1(_03356_),
    .B2(_03357_),
    .X(\u_timer.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__o21a_1 _08009_ (.A1(net1275),
    .A2(\u_timer.u_reg.reg_2[23] ),
    .B1(net1260),
    .X(_03358_));
 sky130_fd_sc_hd__a221o_1 _08010_ (.A1(net1275),
    .A2(\u_timer.u_reg.reg_1[23] ),
    .B1(net1146),
    .B2(\u_timer.u_reg.reg_3[23] ),
    .C1(_03358_),
    .X(_03359_));
 sky130_fd_sc_hd__o21a_1 _08011_ (.A1(net2259),
    .A2(net1227),
    .B1(_03359_),
    .X(\u_timer.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__o21a_1 _08012_ (.A1(net1271),
    .A2(\u_timer.u_reg.reg_2[24] ),
    .B1(net1258),
    .X(_03360_));
 sky130_fd_sc_hd__a22o_1 _08013_ (.A1(net1271),
    .A2(\u_timer.u_reg.reg_1[24] ),
    .B1(net1143),
    .B2(\u_timer.u_reg.reg_3[24] ),
    .X(_03361_));
 sky130_fd_sc_hd__o22a_1 _08014_ (.A1(\u_timer.u_reg.reg_0[24] ),
    .A2(net1222),
    .B1(_03360_),
    .B2(_03361_),
    .X(\u_timer.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__o21a_1 _08015_ (.A1(net1258),
    .A2(\u_timer.u_reg.reg_1[25] ),
    .B1(net1272),
    .X(_03362_));
 sky130_fd_sc_hd__a22o_1 _08016_ (.A1(net1258),
    .A2(\u_timer.u_reg.reg_2[25] ),
    .B1(net1143),
    .B2(\u_timer.u_reg.reg_3[25] ),
    .X(_03363_));
 sky130_fd_sc_hd__o22a_1 _08017_ (.A1(\u_timer.u_reg.reg_0[25] ),
    .A2(net1222),
    .B1(_03362_),
    .B2(_03363_),
    .X(\u_timer.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__o21a_1 _08018_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_2[26] ),
    .B1(net1258),
    .X(_03364_));
 sky130_fd_sc_hd__a22o_1 _08019_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_1[26] ),
    .B1(net1145),
    .B2(\u_timer.u_reg.reg_3[26] ),
    .X(_03365_));
 sky130_fd_sc_hd__o22a_1 _08020_ (.A1(\u_timer.u_reg.reg_0[26] ),
    .A2(net1222),
    .B1(_03364_),
    .B2(_03365_),
    .X(\u_timer.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__o21a_1 _08021_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_2[27] ),
    .B1(net1260),
    .X(_03366_));
 sky130_fd_sc_hd__a221o_1 _08022_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_1[27] ),
    .B1(net1145),
    .B2(\u_timer.u_reg.reg_3[27] ),
    .C1(_03366_),
    .X(_03367_));
 sky130_fd_sc_hd__o21a_1 _08023_ (.A1(net2344),
    .A2(net1228),
    .B1(_03367_),
    .X(\u_timer.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__o21a_1 _08024_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_2[28] ),
    .B1(net1258),
    .X(_03368_));
 sky130_fd_sc_hd__a221o_1 _08025_ (.A1(net1277),
    .A2(\u_timer.u_reg.reg_1[28] ),
    .B1(net1145),
    .B2(\u_timer.u_reg.reg_3[28] ),
    .C1(_03368_),
    .X(_03369_));
 sky130_fd_sc_hd__o21a_1 _08026_ (.A1(net2333),
    .A2(net1228),
    .B1(_03369_),
    .X(\u_timer.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__o21a_1 _08027_ (.A1(net1272),
    .A2(\u_timer.u_reg.reg_2[29] ),
    .B1(net1258),
    .X(_03370_));
 sky130_fd_sc_hd__a221o_1 _08028_ (.A1(net1271),
    .A2(\u_timer.u_reg.reg_1[29] ),
    .B1(net1143),
    .B2(\u_timer.u_reg.reg_3[29] ),
    .C1(_03370_),
    .X(_03371_));
 sky130_fd_sc_hd__o21a_1 _08029_ (.A1(net2320),
    .A2(net1225),
    .B1(_03371_),
    .X(\u_timer.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__o21a_1 _08030_ (.A1(net1272),
    .A2(\u_timer.u_reg.reg_2[30] ),
    .B1(net1258),
    .X(_03372_));
 sky130_fd_sc_hd__a221o_1 _08031_ (.A1(net1271),
    .A2(\u_timer.u_reg.reg_1[30] ),
    .B1(net1143),
    .B2(\u_timer.u_reg.reg_3[30] ),
    .C1(_03372_),
    .X(_03373_));
 sky130_fd_sc_hd__o21a_1 _08032_ (.A1(net2331),
    .A2(net1222),
    .B1(_03373_),
    .X(\u_timer.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__o21a_1 _08033_ (.A1(net1272),
    .A2(\u_timer.u_reg.reg_2[31] ),
    .B1(net1258),
    .X(_03374_));
 sky130_fd_sc_hd__a221o_1 _08034_ (.A1(net1272),
    .A2(\u_timer.u_reg.reg_1[31] ),
    .B1(net1143),
    .B2(\u_timer.u_reg.reg_3[31] ),
    .C1(_03374_),
    .X(_03375_));
 sky130_fd_sc_hd__o21a_1 _08035_ (.A1(\u_timer.u_reg.reg_0[31] ),
    .A2(net1222),
    .B1(_03375_),
    .X(\u_timer.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__mux2_1 _08036_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][0] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][0] ),
    .S(net1080),
    .X(_03376_));
 sky130_fd_sc_hd__mux2_1 _08037_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][0] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][0] ),
    .S(net1084),
    .X(_03377_));
 sky130_fd_sc_hd__a22o_1 _08038_ (.A1(\u_ws281x.u_reg.gfifo[0].u_fifo.full ),
    .A2(net1140),
    .B1(net1135),
    .B2(\u_ws281x.port0_enb ),
    .X(_03378_));
 sky130_fd_sc_hd__a22o_1 _08039_ (.A1(net710),
    .A2(_03376_),
    .B1(_03377_),
    .B2(net714),
    .X(_03379_));
 sky130_fd_sc_hd__a221o_1 _08040_ (.A1(\u_ws281x.cfg_reset_period[0] ),
    .A2(net706),
    .B1(net696),
    .B2(\u_ws281x.cfg_clk_period[0] ),
    .C1(_03378_),
    .X(_03380_));
 sky130_fd_sc_hd__or2_1 _08041_ (.A(_03379_),
    .B(_03380_),
    .X(\u_ws281x.u_reg.reg_out[0] ));
 sky130_fd_sc_hd__mux2_1 _08042_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][1] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][1] ),
    .S(net1080),
    .X(_03381_));
 sky130_fd_sc_hd__mux2_2 _08043_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][1] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][1] ),
    .S(net1084),
    .X(_03382_));
 sky130_fd_sc_hd__a22o_1 _08044_ (.A1(net708),
    .A2(_03381_),
    .B1(_03382_),
    .B2(net714),
    .X(_03383_));
 sky130_fd_sc_hd__a22o_1 _08045_ (.A1(\u_ws281x.cfg_reset_period[1] ),
    .A2(net706),
    .B1(net1135),
    .B2(net2329),
    .X(_03384_));
 sky130_fd_sc_hd__a22o_1 _08046_ (.A1(\u_ws281x.cfg_clk_period[1] ),
    .A2(net696),
    .B1(net1140),
    .B2(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .X(_03385_));
 sky130_fd_sc_hd__or3_1 _08047_ (.A(_03383_),
    .B(_03384_),
    .C(_03385_),
    .X(\u_ws281x.u_reg.reg_out[1] ));
 sky130_fd_sc_hd__a22o_1 _08048_ (.A1(\u_ws281x.cfg_clk_period[2] ),
    .A2(net696),
    .B1(net1135),
    .B2(net2144),
    .X(_03386_));
 sky130_fd_sc_hd__mux2_1 _08049_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][2] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][2] ),
    .S(net1082),
    .X(_03387_));
 sky130_fd_sc_hd__mux2_1 _08050_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][2] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][2] ),
    .S(net1084),
    .X(_03388_));
 sky130_fd_sc_hd__a22o_1 _08051_ (.A1(net708),
    .A2(_03387_),
    .B1(_03388_),
    .B2(net712),
    .X(_03389_));
 sky130_fd_sc_hd__a211o_1 _08052_ (.A1(\u_ws281x.cfg_reset_period[2] ),
    .A2(net705),
    .B1(_03386_),
    .C1(_03389_),
    .X(\u_ws281x.u_reg.reg_out[2] ));
 sky130_fd_sc_hd__a22o_1 _08053_ (.A1(\u_ws281x.cfg_reset_period[3] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_clk_period[3] ),
    .X(_03390_));
 sky130_fd_sc_hd__mux2_1 _08054_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][3] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][3] ),
    .S(net1081),
    .X(_03391_));
 sky130_fd_sc_hd__mux2_1 _08055_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][3] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][3] ),
    .S(net1084),
    .X(_03392_));
 sky130_fd_sc_hd__a22o_1 _08056_ (.A1(net710),
    .A2(_03391_),
    .B1(_03392_),
    .B2(net712),
    .X(_03393_));
 sky130_fd_sc_hd__a211o_1 _08057_ (.A1(net2006),
    .A2(net1135),
    .B1(_03390_),
    .C1(_03393_),
    .X(\u_ws281x.u_reg.reg_out[3] ));
 sky130_fd_sc_hd__a22o_1 _08058_ (.A1(\u_ws281x.cfg_reset_period[4] ),
    .A2(net706),
    .B1(net1140),
    .B2(net2302),
    .X(_03394_));
 sky130_fd_sc_hd__mux2_1 _08059_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][4] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][4] ),
    .S(net1082),
    .X(_03395_));
 sky130_fd_sc_hd__mux2_1 _08060_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][4] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][4] ),
    .S(net1084),
    .X(_03396_));
 sky130_fd_sc_hd__a22o_1 _08061_ (.A1(net708),
    .A2(_03395_),
    .B1(_03396_),
    .B2(net712),
    .X(_03397_));
 sky130_fd_sc_hd__a211o_1 _08062_ (.A1(\u_ws281x.cfg_clk_period[4] ),
    .A2(net695),
    .B1(_03394_),
    .C1(_03397_),
    .X(\u_ws281x.u_reg.reg_out[4] ));
 sky130_fd_sc_hd__a22o_1 _08063_ (.A1(\u_ws281x.cfg_clk_period[5] ),
    .A2(net695),
    .B1(net1140),
    .B2(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .X(_03398_));
 sky130_fd_sc_hd__mux2_1 _08064_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][5] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][5] ),
    .S(net1082),
    .X(_03399_));
 sky130_fd_sc_hd__mux2_1 _08065_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][5] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][5] ),
    .S(net1084),
    .X(_03400_));
 sky130_fd_sc_hd__a22o_1 _08066_ (.A1(net708),
    .A2(_03399_),
    .B1(_03400_),
    .B2(net712),
    .X(_03401_));
 sky130_fd_sc_hd__a211o_1 _08067_ (.A1(\u_ws281x.cfg_reset_period[5] ),
    .A2(net705),
    .B1(_03398_),
    .C1(_03401_),
    .X(\u_ws281x.u_reg.reg_out[5] ));
 sky130_fd_sc_hd__mux2_1 _08068_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][6] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][6] ),
    .S(net1085),
    .X(_03402_));
 sky130_fd_sc_hd__mux2_1 _08069_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][6] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][6] ),
    .S(net1081),
    .X(_03403_));
 sky130_fd_sc_hd__a22o_1 _08070_ (.A1(net712),
    .A2(_03402_),
    .B1(_03403_),
    .B2(net710),
    .X(_03404_));
 sky130_fd_sc_hd__a221o_1 _08071_ (.A1(\u_ws281x.cfg_reset_period[6] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_clk_period[6] ),
    .C1(_03404_),
    .X(\u_ws281x.u_reg.reg_out[6] ));
 sky130_fd_sc_hd__mux2_1 _08072_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][7] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][7] ),
    .S(net1085),
    .X(_03405_));
 sky130_fd_sc_hd__mux2_1 _08073_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][7] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][7] ),
    .S(net1082),
    .X(_03406_));
 sky130_fd_sc_hd__a22o_1 _08074_ (.A1(net712),
    .A2(_03405_),
    .B1(_03406_),
    .B2(net708),
    .X(_03407_));
 sky130_fd_sc_hd__a221o_1 _08075_ (.A1(\u_ws281x.cfg_reset_period[7] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_clk_period[7] ),
    .C1(_03407_),
    .X(\u_ws281x.u_reg.reg_out[7] ));
 sky130_fd_sc_hd__mux2_1 _08076_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][8] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][8] ),
    .S(net1082),
    .X(_03408_));
 sky130_fd_sc_hd__mux2_1 _08077_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][8] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][8] ),
    .S(net1085),
    .X(_03409_));
 sky130_fd_sc_hd__a22o_1 _08078_ (.A1(net708),
    .A2(_03408_),
    .B1(_03409_),
    .B2(net712),
    .X(_03410_));
 sky130_fd_sc_hd__a221o_1 _08079_ (.A1(\u_ws281x.cfg_reset_period[8] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_clk_period[8] ),
    .C1(_03410_),
    .X(\u_ws281x.u_reg.reg_out[8] ));
 sky130_fd_sc_hd__mux2_1 _08080_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][9] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][9] ),
    .S(net1080),
    .X(_03411_));
 sky130_fd_sc_hd__mux2_1 _08081_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][9] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][9] ),
    .S(net1084),
    .X(_03412_));
 sky130_fd_sc_hd__a22o_1 _08082_ (.A1(net708),
    .A2(_03411_),
    .B1(_03412_),
    .B2(net712),
    .X(_03413_));
 sky130_fd_sc_hd__a221o_1 _08083_ (.A1(\u_ws281x.cfg_reset_period[9] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_clk_period[9] ),
    .C1(_03413_),
    .X(\u_ws281x.u_reg.reg_out[9] ));
 sky130_fd_sc_hd__mux2_1 _08084_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][10] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][10] ),
    .S(net1082),
    .X(_03414_));
 sky130_fd_sc_hd__mux2_1 _08085_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][10] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][10] ),
    .S(net1084),
    .X(_03415_));
 sky130_fd_sc_hd__a22o_1 _08086_ (.A1(net708),
    .A2(_03414_),
    .B1(_03415_),
    .B2(net714),
    .X(_03416_));
 sky130_fd_sc_hd__a221o_1 _08087_ (.A1(\u_ws281x.cfg_reset_period[10] ),
    .A2(net705),
    .B1(net696),
    .B2(\u_ws281x.cfg_th0_period[0] ),
    .C1(_03416_),
    .X(\u_ws281x.u_reg.reg_out[10] ));
 sky130_fd_sc_hd__mux2_1 _08088_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][11] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][11] ),
    .S(net1085),
    .X(_03417_));
 sky130_fd_sc_hd__mux2_1 _08089_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][11] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][11] ),
    .S(net1081),
    .X(_03418_));
 sky130_fd_sc_hd__a22o_1 _08090_ (.A1(net712),
    .A2(_03417_),
    .B1(_03418_),
    .B2(net708),
    .X(_03419_));
 sky130_fd_sc_hd__a221o_1 _08091_ (.A1(\u_ws281x.cfg_reset_period[11] ),
    .A2(net705),
    .B1(net695),
    .B2(\u_ws281x.cfg_th0_period[1] ),
    .C1(_03419_),
    .X(\u_ws281x.u_reg.reg_out[11] ));
 sky130_fd_sc_hd__mux2_1 _08092_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][12] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][12] ),
    .S(net1083),
    .X(_03420_));
 sky130_fd_sc_hd__mux2_1 _08093_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][12] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][12] ),
    .S(net1081),
    .X(_03421_));
 sky130_fd_sc_hd__a22o_1 _08094_ (.A1(net712),
    .A2(_03420_),
    .B1(_03421_),
    .B2(net708),
    .X(_03422_));
 sky130_fd_sc_hd__a221o_1 _08095_ (.A1(net2319),
    .A2(net705),
    .B1(net696),
    .B2(\u_ws281x.cfg_th0_period[2] ),
    .C1(_03422_),
    .X(\u_ws281x.u_reg.reg_out[12] ));
 sky130_fd_sc_hd__mux2_1 _08096_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][13] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][13] ),
    .S(net1083),
    .X(_03423_));
 sky130_fd_sc_hd__mux2_1 _08097_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][13] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][13] ),
    .S(net1081),
    .X(_03424_));
 sky130_fd_sc_hd__a22o_1 _08098_ (.A1(net713),
    .A2(_03423_),
    .B1(_03424_),
    .B2(net709),
    .X(_03425_));
 sky130_fd_sc_hd__a221o_1 _08099_ (.A1(\u_ws281x.cfg_reset_period[13] ),
    .A2(net706),
    .B1(net694),
    .B2(\u_ws281x.cfg_th0_period[3] ),
    .C1(_03425_),
    .X(\u_ws281x.u_reg.reg_out[13] ));
 sky130_fd_sc_hd__mux2_1 _08100_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][14] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][14] ),
    .S(net1081),
    .X(_03426_));
 sky130_fd_sc_hd__mux2_1 _08101_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][14] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][14] ),
    .S(net1083),
    .X(_03427_));
 sky130_fd_sc_hd__a22o_1 _08102_ (.A1(net709),
    .A2(_03426_),
    .B1(_03427_),
    .B2(net713),
    .X(_03428_));
 sky130_fd_sc_hd__a221o_1 _08103_ (.A1(\u_ws281x.cfg_reset_period[14] ),
    .A2(net706),
    .B1(net694),
    .B2(\u_ws281x.cfg_th0_period[4] ),
    .C1(_03428_),
    .X(\u_ws281x.u_reg.reg_out[14] ));
 sky130_fd_sc_hd__mux2_1 _08104_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][15] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][15] ),
    .S(net1081),
    .X(_03429_));
 sky130_fd_sc_hd__mux2_1 _08105_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][15] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][15] ),
    .S(net1083),
    .X(_03430_));
 sky130_fd_sc_hd__a22o_1 _08106_ (.A1(net709),
    .A2(_03429_),
    .B1(_03430_),
    .B2(net713),
    .X(_03431_));
 sky130_fd_sc_hd__a221o_1 _08107_ (.A1(\u_ws281x.cfg_reset_period[15] ),
    .A2(net706),
    .B1(net695),
    .B2(\u_ws281x.cfg_th0_period[5] ),
    .C1(_03431_),
    .X(\u_ws281x.u_reg.reg_out[15] ));
 sky130_fd_sc_hd__mux2_1 _08108_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][16] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][16] ),
    .S(net1085),
    .X(_03432_));
 sky130_fd_sc_hd__mux2_1 _08109_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][16] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][16] ),
    .S(net1081),
    .X(_03433_));
 sky130_fd_sc_hd__a22o_1 _08110_ (.A1(net713),
    .A2(_03432_),
    .B1(_03433_),
    .B2(net709),
    .X(_03434_));
 sky130_fd_sc_hd__a21o_1 _08111_ (.A1(\u_ws281x.cfg_th0_period[6] ),
    .A2(net694),
    .B1(_03434_),
    .X(\u_ws281x.u_reg.reg_out[16] ));
 sky130_fd_sc_hd__mux2_1 _08112_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][17] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][17] ),
    .S(net1085),
    .X(_03435_));
 sky130_fd_sc_hd__mux2_1 _08113_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][17] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][17] ),
    .S(net1081),
    .X(_03436_));
 sky130_fd_sc_hd__a22o_1 _08114_ (.A1(net713),
    .A2(_03435_),
    .B1(_03436_),
    .B2(net709),
    .X(_03437_));
 sky130_fd_sc_hd__a21o_1 _08115_ (.A1(\u_ws281x.cfg_th0_period[7] ),
    .A2(net694),
    .B1(_03437_),
    .X(\u_ws281x.u_reg.reg_out[17] ));
 sky130_fd_sc_hd__mux2_1 _08116_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][18] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][18] ),
    .S(net1080),
    .X(_03438_));
 sky130_fd_sc_hd__and3_1 _08117_ (.A(_00996_),
    .B(net1251),
    .C(_03438_),
    .X(_03439_));
 sky130_fd_sc_hd__mux2_1 _08118_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][18] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][18] ),
    .S(net1083),
    .X(_03440_));
 sky130_fd_sc_hd__a221o_1 _08119_ (.A1(\u_ws281x.cfg_th0_period[8] ),
    .A2(net694),
    .B1(_03440_),
    .B2(net713),
    .C1(_03439_),
    .X(\u_ws281x.u_reg.reg_out[18] ));
 sky130_fd_sc_hd__mux2_1 _08120_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][19] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][19] ),
    .S(net1083),
    .X(_03441_));
 sky130_fd_sc_hd__mux2_1 _08121_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][19] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][19] ),
    .S(net1080),
    .X(_03442_));
 sky130_fd_sc_hd__a22o_1 _08122_ (.A1(net713),
    .A2(_03441_),
    .B1(_03442_),
    .B2(net709),
    .X(_03443_));
 sky130_fd_sc_hd__a21o_1 _08123_ (.A1(\u_ws281x.cfg_th0_period[9] ),
    .A2(net694),
    .B1(_03443_),
    .X(\u_ws281x.u_reg.reg_out[19] ));
 sky130_fd_sc_hd__mux2_1 _08124_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][20] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][20] ),
    .S(net1080),
    .X(_03444_));
 sky130_fd_sc_hd__mux2_1 _08125_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][20] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][20] ),
    .S(net1083),
    .X(_03445_));
 sky130_fd_sc_hd__and3_1 _08126_ (.A(net1182),
    .B(net1180),
    .C(_03445_),
    .X(_03446_));
 sky130_fd_sc_hd__a221o_1 _08127_ (.A1(\u_ws281x.cfg_th1_period[0] ),
    .A2(net694),
    .B1(_03444_),
    .B2(net709),
    .C1(_03446_),
    .X(\u_ws281x.u_reg.reg_out[20] ));
 sky130_fd_sc_hd__mux2_1 _08128_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][21] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][21] ),
    .S(net1083),
    .X(_03447_));
 sky130_fd_sc_hd__mux2_1 _08129_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][21] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][21] ),
    .S(net1080),
    .X(_03448_));
 sky130_fd_sc_hd__a22o_1 _08130_ (.A1(net713),
    .A2(_03447_),
    .B1(_03448_),
    .B2(net709),
    .X(_03449_));
 sky130_fd_sc_hd__a21o_1 _08131_ (.A1(\u_ws281x.cfg_th1_period[1] ),
    .A2(net694),
    .B1(_03449_),
    .X(\u_ws281x.u_reg.reg_out[21] ));
 sky130_fd_sc_hd__mux2_1 _08132_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][22] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][22] ),
    .S(net1080),
    .X(_03450_));
 sky130_fd_sc_hd__mux2_1 _08133_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][22] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][22] ),
    .S(net1083),
    .X(_03451_));
 sky130_fd_sc_hd__and3_1 _08134_ (.A(net1182),
    .B(net1180),
    .C(_03451_),
    .X(_03452_));
 sky130_fd_sc_hd__a221o_1 _08135_ (.A1(\u_ws281x.cfg_th1_period[2] ),
    .A2(net694),
    .B1(_03450_),
    .B2(net709),
    .C1(_03452_),
    .X(\u_ws281x.u_reg.reg_out[22] ));
 sky130_fd_sc_hd__mux2_1 _08136_ (.A0(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][23] ),
    .A1(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][23] ),
    .S(net1083),
    .X(_03453_));
 sky130_fd_sc_hd__mux2_1 _08137_ (.A0(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][23] ),
    .A1(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][23] ),
    .S(net1081),
    .X(_03454_));
 sky130_fd_sc_hd__a22o_1 _08138_ (.A1(net713),
    .A2(_03453_),
    .B1(_03454_),
    .B2(net709),
    .X(_03455_));
 sky130_fd_sc_hd__a21o_1 _08139_ (.A1(\u_ws281x.cfg_th1_period[3] ),
    .A2(net694),
    .B1(_03455_),
    .X(\u_ws281x.u_reg.reg_out[23] ));
 sky130_fd_sc_hd__and3_1 _08140_ (.A(\u_ws281x.cfg_th1_period[4] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[24] ));
 sky130_fd_sc_hd__and3_1 _08141_ (.A(\u_ws281x.cfg_th1_period[5] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[25] ));
 sky130_fd_sc_hd__and3_1 _08142_ (.A(\u_ws281x.cfg_th1_period[6] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[26] ));
 sky130_fd_sc_hd__and3_1 _08143_ (.A(\u_ws281x.cfg_th1_period[7] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[27] ));
 sky130_fd_sc_hd__and3_1 _08144_ (.A(\u_ws281x.cfg_th1_period[8] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[28] ));
 sky130_fd_sc_hd__and3_1 _08145_ (.A(\u_ws281x.cfg_th1_period[9] ),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[29] ));
 sky130_fd_sc_hd__and3_1 _08146_ (.A(net2114),
    .B(net1164),
    .C(_01129_),
    .X(\u_ws281x.u_reg.reg_out[30] ));
 sky130_fd_sc_hd__and3_1 _08147_ (.A(net2112),
    .B(net1164),
    .C(net1216),
    .X(\u_ws281x.u_reg.reg_out[31] ));
 sky130_fd_sc_hd__nor3b_1 _08148_ (.A(\u_pwm.blk_sel[2] ),
    .B(\u_pwm.blk_sel[0] ),
    .C_N(net1210),
    .Y(_03456_));
 sky130_fd_sc_hd__and2b_1 _08149_ (.A_N(\u_pwm.blk_sel[2] ),
    .B(\u_pwm.blk_sel[0] ),
    .X(_03457_));
 sky130_fd_sc_hd__nand2b_2 _08150_ (.A_N(\u_pwm.reg_rdata_pwm2[0] ),
    .B(net1209),
    .Y(_03458_));
 sky130_fd_sc_hd__a22o_1 _08151_ (.A1(\u_pwm.reg_rdata_pwm1[0] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03458_),
    .X(_03459_));
 sky130_fd_sc_hd__or3b_1 _08152_ (.A(\u_pwm.blk_sel[2] ),
    .B(net1210),
    .C_N(\u_pwm.blk_sel[0] ),
    .X(_03460_));
 sky130_fd_sc_hd__or2_1 _08153_ (.A(\u_pwm.reg_rdata_pwm0[0] ),
    .B(net1113),
    .X(_03461_));
 sky130_fd_sc_hd__nor3_4 _08154_ (.A(\u_pwm.blk_sel[2] ),
    .B(\u_pwm.blk_sel[0] ),
    .C(net1210),
    .Y(_03462_));
 sky130_fd_sc_hd__a221o_2 _08155_ (.A1(_03459_),
    .A2(_03461_),
    .B1(net1110),
    .B2(\u_pwm.reg_rdata_glbl[0] ),
    .C1(net1092),
    .X(_03463_));
 sky130_fd_sc_hd__and3b_2 _08156_ (.A_N(net1090),
    .B(_00986_),
    .C(\reg_blk_sel[1] ),
    .X(_03464_));
 sky130_fd_sc_hd__or3b_1 _08157_ (.A(net1090),
    .B(\reg_blk_sel[2] ),
    .C_N(\reg_blk_sel[1] ),
    .X(_03465_));
 sky130_fd_sc_hd__nor2_1 _08158_ (.A(net1091),
    .B(_03465_),
    .Y(_03466_));
 sky130_fd_sc_hd__or2_2 _08159_ (.A(net1091),
    .B(_03465_),
    .X(_03467_));
 sky130_fd_sc_hd__o211a_1 _08160_ (.A1(net723),
    .A2(\u_timer.reg_rdata[0] ),
    .B1(_03463_),
    .C1(net559),
    .X(_03468_));
 sky130_fd_sc_hd__nor2_1 _08161_ (.A(\reg_blk_sel[1] ),
    .B(net1090),
    .Y(_03469_));
 sky130_fd_sc_hd__and3_2 _08162_ (.A(net1091),
    .B(\reg_blk_sel[2] ),
    .C(_03469_),
    .X(_03470_));
 sky130_fd_sc_hd__and3_2 _08163_ (.A(net723),
    .B(\reg_blk_sel[2] ),
    .C(_03469_),
    .X(_03471_));
 sky130_fd_sc_hd__or3b_2 _08164_ (.A(net1091),
    .B(_00986_),
    .C_N(_03469_),
    .X(_03472_));
 sky130_fd_sc_hd__a221o_2 _08165_ (.A1(net1086),
    .A2(net66),
    .B1(\u_ws281x.reg_rdata[0] ),
    .B2(net553),
    .C1(net552),
    .X(_03473_));
 sky130_fd_sc_hd__or2_1 _08166_ (.A(\u_semaphore.reg_rdata[0] ),
    .B(net549),
    .X(_03474_));
 sky130_fd_sc_hd__and3_2 _08167_ (.A(net1091),
    .B(_00986_),
    .C(_03469_),
    .X(_03475_));
 sky130_fd_sc_hd__or3b_4 _08168_ (.A(net724),
    .B(\reg_blk_sel[2] ),
    .C_N(_03469_),
    .X(_03476_));
 sky130_fd_sc_hd__and3_1 _08169_ (.A(net724),
    .B(_00986_),
    .C(_03469_),
    .X(_03477_));
 sky130_fd_sc_hd__or4_1 _08170_ (.A(\reg_blk_sel[1] ),
    .B(net1091),
    .C(net1090),
    .D(\reg_blk_sel[2] ),
    .X(_03478_));
 sky130_fd_sc_hd__a221o_1 _08171_ (.A1(_03473_),
    .A2(_03474_),
    .B1(net546),
    .B2(\u_gpio.reg_rdata[0] ),
    .C1(net542),
    .X(_03479_));
 sky130_fd_sc_hd__o22a_2 _08172_ (.A1(net1744),
    .A2(net584),
    .B1(_03479_),
    .B2(_03468_),
    .X(net418));
 sky130_fd_sc_hd__nand2b_2 _08173_ (.A_N(\u_pwm.reg_rdata_pwm2[1] ),
    .B(net1209),
    .Y(_03480_));
 sky130_fd_sc_hd__a22o_1 _08174_ (.A1(\u_pwm.reg_rdata_pwm1[1] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03480_),
    .X(_03481_));
 sky130_fd_sc_hd__or2_1 _08175_ (.A(\u_pwm.reg_rdata_pwm0[1] ),
    .B(net1113),
    .X(_03482_));
 sky130_fd_sc_hd__a221o_2 _08176_ (.A1(\u_pwm.reg_rdata_glbl[1] ),
    .A2(_03462_),
    .B1(_03481_),
    .B2(_03482_),
    .C1(net1091),
    .X(_03483_));
 sky130_fd_sc_hd__o211a_1 _08177_ (.A1(net723),
    .A2(\u_timer.reg_rdata[1] ),
    .B1(net559),
    .C1(_03483_),
    .X(_03484_));
 sky130_fd_sc_hd__a221o_2 _08178_ (.A1(net1086),
    .A2(net77),
    .B1(\u_ws281x.reg_rdata[1] ),
    .B2(net553),
    .C1(net552),
    .X(_03485_));
 sky130_fd_sc_hd__or2_1 _08179_ (.A(\u_semaphore.reg_rdata[1] ),
    .B(net549),
    .X(_03486_));
 sky130_fd_sc_hd__a221o_1 _08180_ (.A1(\u_gpio.reg_rdata[1] ),
    .A2(net547),
    .B1(_03485_),
    .B2(_03486_),
    .C1(net542),
    .X(_03487_));
 sky130_fd_sc_hd__o22a_2 _08181_ (.A1(net1741),
    .A2(net586),
    .B1(_03484_),
    .B2(_03487_),
    .X(net429));
 sky130_fd_sc_hd__nand2b_2 _08182_ (.A_N(\u_pwm.reg_rdata_pwm2[2] ),
    .B(net1209),
    .Y(_03488_));
 sky130_fd_sc_hd__a22o_1 _08183_ (.A1(\u_pwm.reg_rdata_pwm1[2] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03488_),
    .X(_03489_));
 sky130_fd_sc_hd__or2_1 _08184_ (.A(\u_pwm.reg_rdata_pwm0[2] ),
    .B(net1113),
    .X(_03490_));
 sky130_fd_sc_hd__a221o_2 _08185_ (.A1(\u_pwm.reg_rdata_glbl[2] ),
    .A2(_03462_),
    .B1(_03489_),
    .B2(_03490_),
    .C1(net1091),
    .X(_03491_));
 sky130_fd_sc_hd__o211a_1 _08186_ (.A1(net723),
    .A2(\u_timer.reg_rdata[2] ),
    .B1(net559),
    .C1(_03491_),
    .X(_03492_));
 sky130_fd_sc_hd__a221o_2 _08187_ (.A1(net1086),
    .A2(net88),
    .B1(\u_ws281x.reg_rdata[2] ),
    .B2(net553),
    .C1(net552),
    .X(_03493_));
 sky130_fd_sc_hd__or2_1 _08188_ (.A(\u_semaphore.reg_rdata[2] ),
    .B(net549),
    .X(_03494_));
 sky130_fd_sc_hd__a221o_1 _08189_ (.A1(\u_gpio.reg_rdata[2] ),
    .A2(net546),
    .B1(_03493_),
    .B2(_03494_),
    .C1(net542),
    .X(_03495_));
 sky130_fd_sc_hd__o22a_2 _08190_ (.A1(net1747),
    .A2(net586),
    .B1(_03492_),
    .B2(_03495_),
    .X(net440));
 sky130_fd_sc_hd__nand2b_2 _08191_ (.A_N(\u_pwm.reg_rdata_pwm2[3] ),
    .B(net1209),
    .Y(_03496_));
 sky130_fd_sc_hd__a22o_1 _08192_ (.A1(\u_pwm.reg_rdata_pwm1[3] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03496_),
    .X(_03497_));
 sky130_fd_sc_hd__or2_1 _08193_ (.A(\u_pwm.reg_rdata_pwm0[3] ),
    .B(net1113),
    .X(_03498_));
 sky130_fd_sc_hd__a221o_2 _08194_ (.A1(\u_pwm.reg_rdata_glbl[3] ),
    .A2(_03462_),
    .B1(_03497_),
    .B2(_03498_),
    .C1(net1092),
    .X(_03499_));
 sky130_fd_sc_hd__o211a_1 _08195_ (.A1(net724),
    .A2(\u_timer.reg_rdata[3] ),
    .B1(net559),
    .C1(_03499_),
    .X(_03500_));
 sky130_fd_sc_hd__a221o_2 _08196_ (.A1(net1086),
    .A2(net91),
    .B1(\u_ws281x.reg_rdata[3] ),
    .B2(net553),
    .C1(net552),
    .X(_03501_));
 sky130_fd_sc_hd__or2_1 _08197_ (.A(\u_semaphore.reg_rdata[3] ),
    .B(net549),
    .X(_03502_));
 sky130_fd_sc_hd__a221o_1 _08198_ (.A1(\u_gpio.reg_rdata[3] ),
    .A2(net547),
    .B1(_03501_),
    .B2(_03502_),
    .C1(net542),
    .X(_03503_));
 sky130_fd_sc_hd__o22a_2 _08199_ (.A1(net1750),
    .A2(net585),
    .B1(_03500_),
    .B2(_03503_),
    .X(net443));
 sky130_fd_sc_hd__nand2b_2 _08200_ (.A_N(\u_pwm.reg_rdata_pwm2[4] ),
    .B(net1209),
    .Y(_03504_));
 sky130_fd_sc_hd__a22o_1 _08201_ (.A1(\u_pwm.reg_rdata_pwm1[4] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03504_),
    .X(_03505_));
 sky130_fd_sc_hd__or2_1 _08202_ (.A(\u_pwm.reg_rdata_pwm0[4] ),
    .B(net1113),
    .X(_03506_));
 sky130_fd_sc_hd__a221o_2 _08203_ (.A1(\u_pwm.reg_rdata_glbl[4] ),
    .A2(net1110),
    .B1(_03505_),
    .B2(_03506_),
    .C1(net1092),
    .X(_03507_));
 sky130_fd_sc_hd__o211a_1 _08204_ (.A1(net723),
    .A2(\u_timer.reg_rdata[4] ),
    .B1(net559),
    .C1(_03507_),
    .X(_03508_));
 sky130_fd_sc_hd__a221o_2 _08205_ (.A1(net1086),
    .A2(net92),
    .B1(\u_ws281x.reg_rdata[4] ),
    .B2(net554),
    .C1(net551),
    .X(_03509_));
 sky130_fd_sc_hd__or2_1 _08206_ (.A(\u_semaphore.reg_rdata[4] ),
    .B(net549),
    .X(_03510_));
 sky130_fd_sc_hd__a221o_1 _08207_ (.A1(\u_gpio.reg_rdata[4] ),
    .A2(net546),
    .B1(_03509_),
    .B2(_03510_),
    .C1(net542),
    .X(_03511_));
 sky130_fd_sc_hd__o22a_2 _08208_ (.A1(net1753),
    .A2(net584),
    .B1(_03508_),
    .B2(_03511_),
    .X(net444));
 sky130_fd_sc_hd__nand2b_2 _08209_ (.A_N(\u_pwm.reg_rdata_pwm2[5] ),
    .B(net1209),
    .Y(_03512_));
 sky130_fd_sc_hd__a22o_1 _08210_ (.A1(\u_pwm.reg_rdata_pwm1[5] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03512_),
    .X(_03513_));
 sky130_fd_sc_hd__or2_1 _08211_ (.A(\u_pwm.reg_rdata_pwm0[5] ),
    .B(net1113),
    .X(_03514_));
 sky130_fd_sc_hd__a221o_2 _08212_ (.A1(\u_pwm.reg_rdata_glbl[5] ),
    .A2(net1110),
    .B1(_03513_),
    .B2(_03514_),
    .C1(net1092),
    .X(_03515_));
 sky130_fd_sc_hd__o211a_1 _08213_ (.A1(net723),
    .A2(\u_timer.reg_rdata[5] ),
    .B1(net559),
    .C1(_03515_),
    .X(_03516_));
 sky130_fd_sc_hd__a221o_2 _08214_ (.A1(net1087),
    .A2(net93),
    .B1(\u_ws281x.reg_rdata[5] ),
    .B2(net554),
    .C1(net551),
    .X(_03517_));
 sky130_fd_sc_hd__or2_1 _08215_ (.A(\u_semaphore.reg_rdata[5] ),
    .B(net549),
    .X(_03518_));
 sky130_fd_sc_hd__a221o_1 _08216_ (.A1(\u_gpio.reg_rdata[5] ),
    .A2(net546),
    .B1(_03517_),
    .B2(_03518_),
    .C1(net542),
    .X(_03519_));
 sky130_fd_sc_hd__o22a_2 _08217_ (.A1(net1756),
    .A2(net584),
    .B1(_03516_),
    .B2(_03519_),
    .X(net445));
 sky130_fd_sc_hd__a221o_1 _08218_ (.A1(net1087),
    .A2(net94),
    .B1(\u_ws281x.reg_rdata[6] ),
    .B2(net553),
    .C1(net551),
    .X(_03520_));
 sky130_fd_sc_hd__or2_1 _08219_ (.A(\u_semaphore.reg_rdata[6] ),
    .B(net549),
    .X(_03521_));
 sky130_fd_sc_hd__mux2_1 _08220_ (.A0(\u_pwm.reg_rdata_pwm0[6] ),
    .A1(\u_pwm.reg_rdata_pwm2[6] ),
    .S(net1210),
    .X(_03522_));
 sky130_fd_sc_hd__a22o_1 _08221_ (.A1(\u_pwm.reg_rdata_pwm1[6] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03522_),
    .X(_03523_));
 sky130_fd_sc_hd__nor2_1 _08222_ (.A(net724),
    .B(_03465_),
    .Y(_03524_));
 sky130_fd_sc_hd__or2_1 _08223_ (.A(net724),
    .B(_03465_),
    .X(_03525_));
 sky130_fd_sc_hd__a221o_2 _08224_ (.A1(_03520_),
    .A2(_03521_),
    .B1(net540),
    .B2(\u_timer.reg_rdata[6] ),
    .C1(net548),
    .X(_03526_));
 sky130_fd_sc_hd__a21o_1 _08225_ (.A1(net557),
    .A2(_03523_),
    .B1(_03526_),
    .X(_03527_));
 sky130_fd_sc_hd__or2_1 _08226_ (.A(\u_gpio.reg_rdata[6] ),
    .B(_03476_),
    .X(_03528_));
 sky130_fd_sc_hd__a22o_1 _08227_ (.A1(net1735),
    .A2(net541),
    .B1(_03527_),
    .B2(_03528_),
    .X(net446));
 sky130_fd_sc_hd__a221o_1 _08228_ (.A1(net1086),
    .A2(net95),
    .B1(\u_ws281x.reg_rdata[7] ),
    .B2(net554),
    .C1(net552),
    .X(_03529_));
 sky130_fd_sc_hd__or2_1 _08229_ (.A(\u_semaphore.reg_rdata[7] ),
    .B(net550),
    .X(_03530_));
 sky130_fd_sc_hd__mux2_1 _08230_ (.A0(\u_pwm.reg_rdata_pwm0[7] ),
    .A1(\u_pwm.reg_rdata_pwm2[7] ),
    .S(net1729),
    .X(_03531_));
 sky130_fd_sc_hd__a22o_1 _08231_ (.A1(\u_pwm.reg_rdata_pwm1[7] ),
    .A2(net1121),
    .B1(net1116),
    .B2(net1730),
    .X(_03532_));
 sky130_fd_sc_hd__a221o_2 _08232_ (.A1(\u_timer.reg_rdata[7] ),
    .A2(net540),
    .B1(_03529_),
    .B2(_03530_),
    .C1(net548),
    .X(_03533_));
 sky130_fd_sc_hd__a21o_1 _08233_ (.A1(net557),
    .A2(net1731),
    .B1(_03533_),
    .X(_03534_));
 sky130_fd_sc_hd__or2_1 _08234_ (.A(\u_gpio.reg_rdata[7] ),
    .B(_03476_),
    .X(_03535_));
 sky130_fd_sc_hd__a22o_1 _08235_ (.A1(\u_glbl_reg.reg_rdata[7] ),
    .A2(net541),
    .B1(net1732),
    .B2(_03535_),
    .X(net447));
 sky130_fd_sc_hd__nand2b_2 _08236_ (.A_N(\u_pwm.reg_rdata_pwm2[8] ),
    .B(net1207),
    .Y(_03536_));
 sky130_fd_sc_hd__a22o_1 _08237_ (.A1(\u_pwm.reg_rdata_pwm1[8] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03536_),
    .X(_03537_));
 sky130_fd_sc_hd__or2_1 _08238_ (.A(\u_pwm.reg_rdata_pwm0[8] ),
    .B(net1113),
    .X(_03538_));
 sky130_fd_sc_hd__a221o_2 _08239_ (.A1(\u_pwm.reg_rdata_glbl[8] ),
    .A2(net1110),
    .B1(_03537_),
    .B2(_03538_),
    .C1(net1092),
    .X(_03539_));
 sky130_fd_sc_hd__o211a_1 _08240_ (.A1(net723),
    .A2(\u_timer.reg_rdata[8] ),
    .B1(net559),
    .C1(_03539_),
    .X(_03540_));
 sky130_fd_sc_hd__a221o_4 _08241_ (.A1(net1088),
    .A2(net96),
    .B1(\u_ws281x.reg_rdata[8] ),
    .B2(net555),
    .C1(net551),
    .X(_03541_));
 sky130_fd_sc_hd__or2_1 _08242_ (.A(\u_semaphore.reg_rdata[8] ),
    .B(net549),
    .X(_03542_));
 sky130_fd_sc_hd__a221o_1 _08243_ (.A1(\u_gpio.reg_rdata[8] ),
    .A2(net546),
    .B1(_03541_),
    .B2(_03542_),
    .C1(net542),
    .X(_03543_));
 sky130_fd_sc_hd__o22a_2 _08244_ (.A1(net1768),
    .A2(net584),
    .B1(_03540_),
    .B2(_03543_),
    .X(net448));
 sky130_fd_sc_hd__nand2b_2 _08245_ (.A_N(\u_pwm.reg_rdata_pwm2[9] ),
    .B(net1207),
    .Y(_03544_));
 sky130_fd_sc_hd__a22o_1 _08246_ (.A1(\u_pwm.reg_rdata_pwm1[9] ),
    .A2(net1121),
    .B1(net1116),
    .B2(_03544_),
    .X(_03545_));
 sky130_fd_sc_hd__or2_1 _08247_ (.A(\u_pwm.reg_rdata_pwm0[9] ),
    .B(net1112),
    .X(_03546_));
 sky130_fd_sc_hd__a221o_2 _08248_ (.A1(\u_pwm.reg_rdata_glbl[9] ),
    .A2(net1110),
    .B1(_03545_),
    .B2(_03546_),
    .C1(net1092),
    .X(_03547_));
 sky130_fd_sc_hd__o211a_1 _08249_ (.A1(net723),
    .A2(\u_timer.reg_rdata[9] ),
    .B1(net559),
    .C1(_03547_),
    .X(_03548_));
 sky130_fd_sc_hd__a221o_2 _08250_ (.A1(net1087),
    .A2(net97),
    .B1(\u_ws281x.reg_rdata[9] ),
    .B2(net555),
    .C1(net552),
    .X(_03549_));
 sky130_fd_sc_hd__or2_1 _08251_ (.A(\u_semaphore.reg_rdata[9] ),
    .B(net549),
    .X(_03550_));
 sky130_fd_sc_hd__a221o_1 _08252_ (.A1(\u_gpio.reg_rdata[9] ),
    .A2(net548),
    .B1(_03549_),
    .B2(_03550_),
    .C1(net543),
    .X(_03551_));
 sky130_fd_sc_hd__o22a_2 _08253_ (.A1(net1759),
    .A2(net584),
    .B1(_03548_),
    .B2(_03551_),
    .X(net449));
 sky130_fd_sc_hd__nand2b_2 _08254_ (.A_N(\u_pwm.reg_rdata_pwm2[10] ),
    .B(net1729),
    .Y(_03552_));
 sky130_fd_sc_hd__a22o_1 _08255_ (.A1(\u_pwm.reg_rdata_pwm1[10] ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03552_),
    .X(_03553_));
 sky130_fd_sc_hd__or2_1 _08256_ (.A(\u_pwm.reg_rdata_pwm0[10] ),
    .B(net1113),
    .X(_03554_));
 sky130_fd_sc_hd__a221o_1 _08257_ (.A1(\u_pwm.reg_rdata_glbl[10] ),
    .A2(net1110),
    .B1(_03553_),
    .B2(_03554_),
    .C1(net1092),
    .X(_03555_));
 sky130_fd_sc_hd__o211a_1 _08258_ (.A1(net723),
    .A2(\u_timer.reg_rdata[10] ),
    .B1(net559),
    .C1(_03555_),
    .X(_03556_));
 sky130_fd_sc_hd__a221o_2 _08259_ (.A1(net1087),
    .A2(net67),
    .B1(\u_ws281x.reg_rdata[10] ),
    .B2(net553),
    .C1(net551),
    .X(_03557_));
 sky130_fd_sc_hd__or2_1 _08260_ (.A(\u_semaphore.reg_rdata[10] ),
    .B(net549),
    .X(_03558_));
 sky130_fd_sc_hd__a221o_1 _08261_ (.A1(\u_gpio.reg_rdata[10] ),
    .A2(net546),
    .B1(_03557_),
    .B2(_03558_),
    .C1(net542),
    .X(_03559_));
 sky130_fd_sc_hd__o22a_2 _08262_ (.A1(net1762),
    .A2(net584),
    .B1(_03556_),
    .B2(_03559_),
    .X(net419));
 sky130_fd_sc_hd__a221o_1 _08263_ (.A1(net1088),
    .A2(net68),
    .B1(\u_ws281x.reg_rdata[11] ),
    .B2(net555),
    .C1(net551),
    .X(_03560_));
 sky130_fd_sc_hd__or2_1 _08264_ (.A(\u_semaphore.reg_rdata[11] ),
    .B(net550),
    .X(_03561_));
 sky130_fd_sc_hd__mux2_1 _08265_ (.A0(\u_pwm.reg_rdata_pwm0[11] ),
    .A1(\u_pwm.reg_rdata_pwm2[11] ),
    .S(net1210),
    .X(_03562_));
 sky130_fd_sc_hd__a22o_1 _08266_ (.A1(\u_pwm.reg_rdata_pwm1[11] ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03562_),
    .X(_03563_));
 sky130_fd_sc_hd__a221o_2 _08267_ (.A1(\u_timer.reg_rdata[11] ),
    .A2(net540),
    .B1(_03560_),
    .B2(_03561_),
    .C1(net548),
    .X(_03564_));
 sky130_fd_sc_hd__a21o_1 _08268_ (.A1(net557),
    .A2(_03563_),
    .B1(_03564_),
    .X(_03565_));
 sky130_fd_sc_hd__or2_1 _08269_ (.A(\u_gpio.reg_rdata[11] ),
    .B(_03476_),
    .X(_03566_));
 sky130_fd_sc_hd__a22o_1 _08270_ (.A1(net1723),
    .A2(net541),
    .B1(_03565_),
    .B2(_03566_),
    .X(net420));
 sky130_fd_sc_hd__a221o_1 _08271_ (.A1(net1086),
    .A2(net69),
    .B1(\u_ws281x.reg_rdata[12] ),
    .B2(net555),
    .C1(net551),
    .X(_03567_));
 sky130_fd_sc_hd__or2_1 _08272_ (.A(\u_semaphore.reg_rdata[12] ),
    .B(net550),
    .X(_03568_));
 sky130_fd_sc_hd__mux2_1 _08273_ (.A0(\u_pwm.reg_rdata_pwm0[12] ),
    .A1(\u_pwm.reg_rdata_pwm2[12] ),
    .S(net1210),
    .X(_03569_));
 sky130_fd_sc_hd__a22o_1 _08274_ (.A1(\u_pwm.reg_rdata_pwm1[12] ),
    .A2(net1120),
    .B1(net1115),
    .B2(_03569_),
    .X(_03570_));
 sky130_fd_sc_hd__a221o_2 _08275_ (.A1(\u_timer.reg_rdata[12] ),
    .A2(net540),
    .B1(_03567_),
    .B2(_03568_),
    .C1(_03475_),
    .X(_03571_));
 sky130_fd_sc_hd__a21o_1 _08276_ (.A1(net557),
    .A2(_03570_),
    .B1(_03571_),
    .X(_03572_));
 sky130_fd_sc_hd__or2_1 _08277_ (.A(\u_gpio.reg_rdata[12] ),
    .B(_03476_),
    .X(_03573_));
 sky130_fd_sc_hd__a22o_1 _08278_ (.A1(net1717),
    .A2(net541),
    .B1(_03572_),
    .B2(_03573_),
    .X(net421));
 sky130_fd_sc_hd__a221o_1 _08279_ (.A1(net1088),
    .A2(net70),
    .B1(\u_ws281x.reg_rdata[13] ),
    .B2(net555),
    .C1(net551),
    .X(_03574_));
 sky130_fd_sc_hd__or2_1 _08280_ (.A(\u_semaphore.reg_rdata[13] ),
    .B(net550),
    .X(_03575_));
 sky130_fd_sc_hd__mux2_1 _08281_ (.A0(\u_pwm.reg_rdata_pwm0[13] ),
    .A1(\u_pwm.reg_rdata_pwm2[13] ),
    .S(net1210),
    .X(_03576_));
 sky130_fd_sc_hd__a22o_1 _08282_ (.A1(\u_pwm.reg_rdata_pwm1[13] ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03576_),
    .X(_03577_));
 sky130_fd_sc_hd__a221o_2 _08283_ (.A1(\u_timer.reg_rdata[13] ),
    .A2(net540),
    .B1(_03574_),
    .B2(_03575_),
    .C1(_03475_),
    .X(_03578_));
 sky130_fd_sc_hd__a21o_1 _08284_ (.A1(net557),
    .A2(_03577_),
    .B1(_03578_),
    .X(_03579_));
 sky130_fd_sc_hd__or2_1 _08285_ (.A(\u_gpio.reg_rdata[13] ),
    .B(_03476_),
    .X(_03580_));
 sky130_fd_sc_hd__a22o_1 _08286_ (.A1(net1711),
    .A2(net541),
    .B1(_03579_),
    .B2(_03580_),
    .X(net422));
 sky130_fd_sc_hd__a221o_1 _08287_ (.A1(net1088),
    .A2(net71),
    .B1(\u_ws281x.reg_rdata[14] ),
    .B2(net555),
    .C1(net551),
    .X(_03581_));
 sky130_fd_sc_hd__or2_1 _08288_ (.A(\u_semaphore.reg_rdata[14] ),
    .B(net550),
    .X(_03582_));
 sky130_fd_sc_hd__mux2_1 _08289_ (.A0(\u_pwm.reg_rdata_pwm0[14] ),
    .A1(\u_pwm.reg_rdata_pwm2[14] ),
    .S(net1210),
    .X(_03583_));
 sky130_fd_sc_hd__a22o_1 _08290_ (.A1(\u_pwm.reg_rdata_pwm1[14] ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03583_),
    .X(_03584_));
 sky130_fd_sc_hd__a221o_2 _08291_ (.A1(\u_timer.reg_rdata[14] ),
    .A2(net540),
    .B1(_03581_),
    .B2(_03582_),
    .C1(net548),
    .X(_03585_));
 sky130_fd_sc_hd__a21o_1 _08292_ (.A1(_03466_),
    .A2(_03584_),
    .B1(_03585_),
    .X(_03586_));
 sky130_fd_sc_hd__or2_1 _08293_ (.A(\u_gpio.reg_rdata[14] ),
    .B(_03476_),
    .X(_03587_));
 sky130_fd_sc_hd__a22o_1 _08294_ (.A1(net1738),
    .A2(net541),
    .B1(_03586_),
    .B2(_03587_),
    .X(net423));
 sky130_fd_sc_hd__a221o_1 _08295_ (.A1(net1088),
    .A2(net72),
    .B1(\u_ws281x.reg_rdata[15] ),
    .B2(net555),
    .C1(net551),
    .X(_03588_));
 sky130_fd_sc_hd__or2_1 _08296_ (.A(\u_semaphore.reg_rdata[15] ),
    .B(net550),
    .X(_03589_));
 sky130_fd_sc_hd__mux2_1 _08297_ (.A0(\u_pwm.reg_rdata_pwm0[15] ),
    .A1(\u_pwm.reg_rdata_pwm2[15] ),
    .S(net1210),
    .X(_03590_));
 sky130_fd_sc_hd__a22o_1 _08298_ (.A1(\u_pwm.reg_rdata_pwm1[15] ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03590_),
    .X(_03591_));
 sky130_fd_sc_hd__a221o_2 _08299_ (.A1(\u_timer.reg_rdata[15] ),
    .A2(net540),
    .B1(_03588_),
    .B2(_03589_),
    .C1(net548),
    .X(_03592_));
 sky130_fd_sc_hd__a21o_1 _08300_ (.A1(net557),
    .A2(_03591_),
    .B1(_03592_),
    .X(_03593_));
 sky130_fd_sc_hd__or2_1 _08301_ (.A(\u_gpio.reg_rdata[15] ),
    .B(_03476_),
    .X(_03594_));
 sky130_fd_sc_hd__a22o_1 _08302_ (.A1(net1720),
    .A2(net541),
    .B1(_03593_),
    .B2(_03594_),
    .X(net424));
 sky130_fd_sc_hd__nand2b_1 _08303_ (.A_N(\u_pwm.reg_rdata_pwm2[16] ),
    .B(net1209),
    .Y(_03595_));
 sky130_fd_sc_hd__a22o_2 _08304_ (.A1(\u_pwm.reg_rdata_pwm1[16] ),
    .A2(net1123),
    .B1(net1118),
    .B2(_03595_),
    .X(_03596_));
 sky130_fd_sc_hd__or2_1 _08305_ (.A(\u_pwm.reg_rdata_pwm0[16] ),
    .B(net1112),
    .X(_03597_));
 sky130_fd_sc_hd__a22o_1 _08306_ (.A1(\u_pwm.reg_rdata_glbl[16] ),
    .A2(net1110),
    .B1(_03596_),
    .B2(_03597_),
    .X(_03598_));
 sky130_fd_sc_hd__a221o_2 _08307_ (.A1(net1087),
    .A2(net73),
    .B1(\u_ws281x.reg_rdata[16] ),
    .B2(net554),
    .C1(_03464_),
    .X(_03599_));
 sky130_fd_sc_hd__o221a_1 _08308_ (.A1(\u_timer.reg_rdata[16] ),
    .A2(_03525_),
    .B1(_03598_),
    .B2(_03467_),
    .C1(_03599_),
    .X(_03600_));
 sky130_fd_sc_hd__mux2_1 _08309_ (.A0(\u_gpio.reg_rdata[16] ),
    .A1(_03600_),
    .S(_03476_),
    .X(_03601_));
 sky130_fd_sc_hd__a21o_1 _08310_ (.A1(net1726),
    .A2(net544),
    .B1(_03601_),
    .X(net425));
 sky130_fd_sc_hd__nand2b_1 _08311_ (.A_N(\u_pwm.reg_rdata_pwm2[17] ),
    .B(net1207),
    .Y(_03602_));
 sky130_fd_sc_hd__a22o_2 _08312_ (.A1(\u_pwm.reg_rdata_pwm1[17] ),
    .A2(net1120),
    .B1(net1115),
    .B2(_03602_),
    .X(_03603_));
 sky130_fd_sc_hd__or2_1 _08313_ (.A(\u_pwm.reg_rdata_pwm0[17] ),
    .B(net1112),
    .X(_03604_));
 sky130_fd_sc_hd__a221o_1 _08314_ (.A1(\u_pwm.reg_rdata_glbl[17] ),
    .A2(net1110),
    .B1(_03603_),
    .B2(_03604_),
    .C1(_03467_),
    .X(_03605_));
 sky130_fd_sc_hd__a221o_2 _08315_ (.A1(net1087),
    .A2(net74),
    .B1(\u_ws281x.reg_rdata[17] ),
    .B2(net553),
    .C1(_03464_),
    .X(_03606_));
 sky130_fd_sc_hd__o211a_1 _08316_ (.A1(\u_timer.reg_rdata[17] ),
    .A2(_03525_),
    .B1(_03605_),
    .C1(_03606_),
    .X(_03607_));
 sky130_fd_sc_hd__mux2_1 _08317_ (.A0(\u_gpio.reg_rdata[17] ),
    .A1(_03607_),
    .S(_03476_),
    .X(_03608_));
 sky130_fd_sc_hd__a21o_2 _08318_ (.A1(net1708),
    .A2(net544),
    .B1(_03608_),
    .X(net426));
 sky130_fd_sc_hd__nand2b_1 _08319_ (.A_N(\u_pwm.reg_rdata_pwm2[18] ),
    .B(net1209),
    .Y(_03609_));
 sky130_fd_sc_hd__a22o_2 _08320_ (.A1(\u_pwm.reg_rdata_pwm1[18] ),
    .A2(net1123),
    .B1(net1118),
    .B2(_03609_),
    .X(_03610_));
 sky130_fd_sc_hd__or2_1 _08321_ (.A(\u_pwm.reg_rdata_pwm0[18] ),
    .B(net1112),
    .X(_03611_));
 sky130_fd_sc_hd__a221o_1 _08322_ (.A1(\u_pwm.reg_rdata_glbl[18] ),
    .A2(net1110),
    .B1(_03610_),
    .B2(_03611_),
    .C1(_03467_),
    .X(_03612_));
 sky130_fd_sc_hd__a221o_2 _08323_ (.A1(net1087),
    .A2(net75),
    .B1(\u_ws281x.reg_rdata[18] ),
    .B2(net554),
    .C1(_03464_),
    .X(_03613_));
 sky130_fd_sc_hd__o211a_1 _08324_ (.A1(\u_timer.reg_rdata[18] ),
    .A2(_03525_),
    .B1(_03612_),
    .C1(_03613_),
    .X(_03614_));
 sky130_fd_sc_hd__mux2_1 _08325_ (.A0(\u_gpio.reg_rdata[18] ),
    .A1(_03614_),
    .S(_03476_),
    .X(_03615_));
 sky130_fd_sc_hd__a21o_2 _08326_ (.A1(net1714),
    .A2(net544),
    .B1(_03615_),
    .X(net427));
 sky130_fd_sc_hd__a22o_2 _08327_ (.A1(net1086),
    .A2(net76),
    .B1(net1794),
    .B2(net553),
    .X(_03616_));
 sky130_fd_sc_hd__nand2b_1 _08328_ (.A_N(\u_pwm.reg_rdata_pwm2[19] ),
    .B(net1209),
    .Y(_03617_));
 sky130_fd_sc_hd__a22o_2 _08329_ (.A1(\u_pwm.reg_rdata_pwm1[19] ),
    .A2(net1123),
    .B1(net1118),
    .B2(_03617_),
    .X(_03618_));
 sky130_fd_sc_hd__or2_1 _08330_ (.A(\u_pwm.reg_rdata_pwm0[19] ),
    .B(net1112),
    .X(_03619_));
 sky130_fd_sc_hd__a221o_1 _08331_ (.A1(\u_gpio.reg_rdata[19] ),
    .A2(net548),
    .B1(net540),
    .B2(\u_timer.reg_rdata[19] ),
    .C1(net543),
    .X(_03620_));
 sky130_fd_sc_hd__a31o_1 _08332_ (.A1(net558),
    .A2(_03618_),
    .A3(_03619_),
    .B1(_03620_),
    .X(_03621_));
 sky130_fd_sc_hd__o22a_2 _08333_ (.A1(\u_glbl_reg.reg_rdata[19] ),
    .A2(net584),
    .B1(net1795),
    .B2(_03621_),
    .X(net428));
 sky130_fd_sc_hd__a22o_1 _08334_ (.A1(net1086),
    .A2(net78),
    .B1(\u_ws281x.reg_rdata[20] ),
    .B2(net554),
    .X(_03622_));
 sky130_fd_sc_hd__nand2b_1 _08335_ (.A_N(\u_pwm.reg_rdata_pwm2[20] ),
    .B(net1207),
    .Y(_03623_));
 sky130_fd_sc_hd__a22o_2 _08336_ (.A1(\u_pwm.reg_rdata_pwm1[20] ),
    .A2(net1120),
    .B1(net1115),
    .B2(_03623_),
    .X(_03624_));
 sky130_fd_sc_hd__or2_1 _08337_ (.A(\u_pwm.reg_rdata_pwm0[20] ),
    .B(net1111),
    .X(_03625_));
 sky130_fd_sc_hd__a221o_1 _08338_ (.A1(\u_gpio.reg_rdata[20] ),
    .A2(net548),
    .B1(net540),
    .B2(\u_timer.reg_rdata[20] ),
    .C1(net543),
    .X(_03626_));
 sky130_fd_sc_hd__a31o_1 _08339_ (.A1(net558),
    .A2(_03624_),
    .A3(_03625_),
    .B1(_03626_),
    .X(_03627_));
 sky130_fd_sc_hd__o22a_2 _08340_ (.A1(net1811),
    .A2(net585),
    .B1(_03622_),
    .B2(_03627_),
    .X(net430));
 sky130_fd_sc_hd__a22o_2 _08341_ (.A1(net1088),
    .A2(net79),
    .B1(\u_ws281x.reg_rdata[21] ),
    .B2(net555),
    .X(_03628_));
 sky130_fd_sc_hd__nand2b_1 _08342_ (.A_N(\u_pwm.reg_rdata_pwm2[21] ),
    .B(net1208),
    .Y(_03629_));
 sky130_fd_sc_hd__a22o_2 _08343_ (.A1(\u_pwm.reg_rdata_pwm1[21] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03629_),
    .X(_03630_));
 sky130_fd_sc_hd__or2_1 _08344_ (.A(\u_pwm.reg_rdata_pwm0[21] ),
    .B(net1111),
    .X(_03631_));
 sky130_fd_sc_hd__a221o_1 _08345_ (.A1(\u_gpio.reg_rdata[21] ),
    .A2(net548),
    .B1(net540),
    .B2(\u_timer.reg_rdata[21] ),
    .C1(net543),
    .X(_03632_));
 sky130_fd_sc_hd__a31o_1 _08346_ (.A1(net558),
    .A2(_03630_),
    .A3(_03631_),
    .B1(_03632_),
    .X(_03633_));
 sky130_fd_sc_hd__o22a_2 _08347_ (.A1(net1804),
    .A2(net584),
    .B1(_03628_),
    .B2(_03633_),
    .X(net431));
 sky130_fd_sc_hd__a22o_2 _08348_ (.A1(net1086),
    .A2(net80),
    .B1(net1784),
    .B2(net553),
    .X(_03634_));
 sky130_fd_sc_hd__nand2b_1 _08349_ (.A_N(\u_pwm.reg_rdata_pwm2[22] ),
    .B(net1208),
    .Y(_03635_));
 sky130_fd_sc_hd__a22o_2 _08350_ (.A1(\u_pwm.reg_rdata_pwm1[22] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03635_),
    .X(_03636_));
 sky130_fd_sc_hd__or2_1 _08351_ (.A(\u_pwm.reg_rdata_pwm0[22] ),
    .B(net1111),
    .X(_03637_));
 sky130_fd_sc_hd__a221o_1 _08352_ (.A1(\u_gpio.reg_rdata[22] ),
    .A2(net546),
    .B1(net539),
    .B2(\u_timer.reg_rdata[22] ),
    .C1(net542),
    .X(_03638_));
 sky130_fd_sc_hd__a31o_1 _08353_ (.A1(net558),
    .A2(_03636_),
    .A3(_03637_),
    .B1(_03638_),
    .X(_03639_));
 sky130_fd_sc_hd__o22a_2 _08354_ (.A1(\u_glbl_reg.reg_rdata[22] ),
    .A2(net584),
    .B1(net1785),
    .B2(_03639_),
    .X(net432));
 sky130_fd_sc_hd__a22o_2 _08355_ (.A1(net1088),
    .A2(net81),
    .B1(\u_ws281x.reg_rdata[23] ),
    .B2(net555),
    .X(_03640_));
 sky130_fd_sc_hd__nand2b_1 _08356_ (.A_N(\u_pwm.reg_rdata_pwm2[23] ),
    .B(net1207),
    .Y(_03641_));
 sky130_fd_sc_hd__a22o_2 _08357_ (.A1(\u_pwm.reg_rdata_pwm1[23] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03641_),
    .X(_03642_));
 sky130_fd_sc_hd__or2_1 _08358_ (.A(\u_pwm.reg_rdata_pwm0[23] ),
    .B(net1111),
    .X(_03643_));
 sky130_fd_sc_hd__a221o_1 _08359_ (.A1(\u_gpio.reg_rdata[23] ),
    .A2(net546),
    .B1(net539),
    .B2(\u_timer.reg_rdata[23] ),
    .C1(net543),
    .X(_03644_));
 sky130_fd_sc_hd__a31o_1 _08360_ (.A1(net558),
    .A2(_03642_),
    .A3(_03643_),
    .B1(_03644_),
    .X(_03645_));
 sky130_fd_sc_hd__o22a_2 _08361_ (.A1(net1801),
    .A2(net584),
    .B1(_03640_),
    .B2(_03645_),
    .X(net433));
 sky130_fd_sc_hd__a22o_2 _08362_ (.A1(net1088),
    .A2(net82),
    .B1(\u_ws281x.reg_rdata[24] ),
    .B2(net556),
    .X(_03646_));
 sky130_fd_sc_hd__nand2b_1 _08363_ (.A_N(\u_pwm.reg_rdata_pwm2[24] ),
    .B(net1208),
    .Y(_03647_));
 sky130_fd_sc_hd__a22o_1 _08364_ (.A1(\u_pwm.reg_rdata_pwm1[24] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03647_),
    .X(_03648_));
 sky130_fd_sc_hd__or2_1 _08365_ (.A(\u_pwm.reg_rdata_pwm0[24] ),
    .B(net1111),
    .X(_03649_));
 sky130_fd_sc_hd__a221o_1 _08366_ (.A1(\u_gpio.reg_rdata[24] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[24] ),
    .C1(net541),
    .X(_03650_));
 sky130_fd_sc_hd__a31o_1 _08367_ (.A1(net558),
    .A2(_03648_),
    .A3(_03649_),
    .B1(_03650_),
    .X(_03651_));
 sky130_fd_sc_hd__o22a_2 _08368_ (.A1(net1788),
    .A2(net585),
    .B1(_03646_),
    .B2(_03651_),
    .X(net434));
 sky130_fd_sc_hd__a22o_4 _08369_ (.A1(net1088),
    .A2(net83),
    .B1(net1780),
    .B2(net556),
    .X(_03652_));
 sky130_fd_sc_hd__nand2b_1 _08370_ (.A_N(\u_pwm.reg_rdata_pwm2[25] ),
    .B(net1207),
    .Y(_03653_));
 sky130_fd_sc_hd__a22o_1 _08371_ (.A1(\u_pwm.reg_rdata_pwm1[25] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03653_),
    .X(_03654_));
 sky130_fd_sc_hd__or2_1 _08372_ (.A(\u_pwm.reg_rdata_pwm0[25] ),
    .B(net1112),
    .X(_03655_));
 sky130_fd_sc_hd__a221o_1 _08373_ (.A1(\u_gpio.reg_rdata[25] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[25] ),
    .C1(net545),
    .X(_03656_));
 sky130_fd_sc_hd__a31o_1 _08374_ (.A1(net557),
    .A2(_03654_),
    .A3(_03655_),
    .B1(_03656_),
    .X(_03657_));
 sky130_fd_sc_hd__o22a_2 _08375_ (.A1(\u_glbl_reg.reg_rdata[25] ),
    .A2(net586),
    .B1(net1781),
    .B2(_03657_),
    .X(net435));
 sky130_fd_sc_hd__a22o_2 _08376_ (.A1(net1088),
    .A2(net84),
    .B1(\u_ws281x.reg_rdata[26] ),
    .B2(net555),
    .X(_03658_));
 sky130_fd_sc_hd__nand2b_1 _08377_ (.A_N(\u_pwm.reg_rdata_pwm2[26] ),
    .B(net1207),
    .Y(_03659_));
 sky130_fd_sc_hd__a22o_2 _08378_ (.A1(\u_pwm.reg_rdata_pwm1[26] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03659_),
    .X(_03660_));
 sky130_fd_sc_hd__or2_1 _08379_ (.A(\u_pwm.reg_rdata_pwm0[26] ),
    .B(net1112),
    .X(_03661_));
 sky130_fd_sc_hd__a221o_1 _08380_ (.A1(\u_gpio.reg_rdata[26] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[26] ),
    .C1(net541),
    .X(_03662_));
 sky130_fd_sc_hd__a31o_1 _08381_ (.A1(net558),
    .A2(_03660_),
    .A3(_03661_),
    .B1(_03662_),
    .X(_03663_));
 sky130_fd_sc_hd__o22a_2 _08382_ (.A1(net1798),
    .A2(net585),
    .B1(_03658_),
    .B2(_03663_),
    .X(net436));
 sky130_fd_sc_hd__a22o_2 _08383_ (.A1(net1089),
    .A2(net85),
    .B1(net1807),
    .B2(net556),
    .X(_03664_));
 sky130_fd_sc_hd__nand2b_1 _08384_ (.A_N(\u_pwm.reg_rdata_pwm2[27] ),
    .B(net1207),
    .Y(_03665_));
 sky130_fd_sc_hd__a22o_2 _08385_ (.A1(\u_pwm.reg_rdata_pwm1[27] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03665_),
    .X(_03666_));
 sky130_fd_sc_hd__or2_1 _08386_ (.A(\u_pwm.reg_rdata_pwm0[27] ),
    .B(net1112),
    .X(_03667_));
 sky130_fd_sc_hd__a221o_1 _08387_ (.A1(\u_gpio.reg_rdata[27] ),
    .A2(net546),
    .B1(net539),
    .B2(\u_timer.reg_rdata[27] ),
    .C1(net542),
    .X(_03668_));
 sky130_fd_sc_hd__a31o_1 _08388_ (.A1(net558),
    .A2(_03666_),
    .A3(_03667_),
    .B1(_03668_),
    .X(_03669_));
 sky130_fd_sc_hd__o22a_2 _08389_ (.A1(\u_glbl_reg.reg_rdata[27] ),
    .A2(net585),
    .B1(net1808),
    .B2(_03669_),
    .X(net437));
 sky130_fd_sc_hd__a22o_2 _08390_ (.A1(net1089),
    .A2(net86),
    .B1(\u_ws281x.reg_rdata[28] ),
    .B2(net556),
    .X(_03670_));
 sky130_fd_sc_hd__nand2b_1 _08391_ (.A_N(\u_pwm.reg_rdata_pwm2[28] ),
    .B(net1208),
    .Y(_03671_));
 sky130_fd_sc_hd__a22o_1 _08392_ (.A1(\u_pwm.reg_rdata_pwm1[28] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03671_),
    .X(_03672_));
 sky130_fd_sc_hd__or2_1 _08393_ (.A(\u_pwm.reg_rdata_pwm0[28] ),
    .B(net1111),
    .X(_03673_));
 sky130_fd_sc_hd__a221o_1 _08394_ (.A1(\u_gpio.reg_rdata[28] ),
    .A2(net546),
    .B1(net539),
    .B2(\u_timer.reg_rdata[28] ),
    .C1(net541),
    .X(_03674_));
 sky130_fd_sc_hd__a31o_1 _08395_ (.A1(net558),
    .A2(_03672_),
    .A3(_03673_),
    .B1(_03674_),
    .X(_03675_));
 sky130_fd_sc_hd__o22a_2 _08396_ (.A1(net1791),
    .A2(net585),
    .B1(_03670_),
    .B2(_03675_),
    .X(net438));
 sky130_fd_sc_hd__a22o_4 _08397_ (.A1(net1089),
    .A2(net87),
    .B1(net1776),
    .B2(net556),
    .X(_03676_));
 sky130_fd_sc_hd__nand2b_1 _08398_ (.A_N(\u_pwm.reg_rdata_pwm2[29] ),
    .B(net1207),
    .Y(_03677_));
 sky130_fd_sc_hd__a22o_1 _08399_ (.A1(\u_pwm.reg_rdata_pwm1[29] ),
    .A2(net1119),
    .B1(net1114),
    .B2(_03677_),
    .X(_03678_));
 sky130_fd_sc_hd__or2_1 _08400_ (.A(\u_pwm.reg_rdata_pwm0[29] ),
    .B(net1111),
    .X(_03679_));
 sky130_fd_sc_hd__a221o_1 _08401_ (.A1(\u_gpio.reg_rdata[29] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[29] ),
    .C1(net545),
    .X(_03680_));
 sky130_fd_sc_hd__a31o_1 _08402_ (.A1(net557),
    .A2(_03678_),
    .A3(_03679_),
    .B1(_03680_),
    .X(_03681_));
 sky130_fd_sc_hd__o22a_2 _08403_ (.A1(\u_glbl_reg.reg_rdata[29] ),
    .A2(net586),
    .B1(net1777),
    .B2(_03681_),
    .X(net439));
 sky130_fd_sc_hd__a22o_4 _08404_ (.A1(net1089),
    .A2(net89),
    .B1(\u_ws281x.reg_rdata[30] ),
    .B2(net556),
    .X(_03682_));
 sky130_fd_sc_hd__nand2b_1 _08405_ (.A_N(\u_pwm.reg_rdata_pwm2[30] ),
    .B(net1207),
    .Y(_03683_));
 sky130_fd_sc_hd__a22o_1 _08406_ (.A1(net1771),
    .A2(net1119),
    .B1(net1114),
    .B2(_03683_),
    .X(_03684_));
 sky130_fd_sc_hd__or2_1 _08407_ (.A(\u_pwm.reg_rdata_pwm0[30] ),
    .B(net1111),
    .X(_03685_));
 sky130_fd_sc_hd__a221o_1 _08408_ (.A1(\u_gpio.reg_rdata[30] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[30] ),
    .C1(net545),
    .X(_03686_));
 sky130_fd_sc_hd__a31o_1 _08409_ (.A1(net557),
    .A2(net1772),
    .A3(_03685_),
    .B1(_03686_),
    .X(_03687_));
 sky130_fd_sc_hd__o22a_2 _08410_ (.A1(\u_glbl_reg.reg_rdata[30] ),
    .A2(net586),
    .B1(_03682_),
    .B2(net1773),
    .X(net441));
 sky130_fd_sc_hd__a22o_4 _08411_ (.A1(net1089),
    .A2(net90),
    .B1(\u_ws281x.reg_rdata[31] ),
    .B2(net556),
    .X(_03688_));
 sky130_fd_sc_hd__nand2b_1 _08412_ (.A_N(\u_pwm.reg_rdata_pwm2[31] ),
    .B(net1208),
    .Y(_03689_));
 sky130_fd_sc_hd__a22o_1 _08413_ (.A1(\u_pwm.reg_rdata_pwm1[31] ),
    .A2(net1120),
    .B1(net1115),
    .B2(_03689_),
    .X(_03690_));
 sky130_fd_sc_hd__or2_1 _08414_ (.A(\u_pwm.reg_rdata_pwm0[31] ),
    .B(net1111),
    .X(_03691_));
 sky130_fd_sc_hd__a221o_1 _08415_ (.A1(\u_gpio.reg_rdata[31] ),
    .A2(net547),
    .B1(net539),
    .B2(\u_timer.reg_rdata[31] ),
    .C1(net545),
    .X(_03692_));
 sky130_fd_sc_hd__a31o_1 _08416_ (.A1(net557),
    .A2(_03690_),
    .A3(_03691_),
    .B1(_03692_),
    .X(_03693_));
 sky130_fd_sc_hd__o22a_2 _08417_ (.A1(net1765),
    .A2(net586),
    .B1(_03688_),
    .B2(_03693_),
    .X(net442));
 sky130_fd_sc_hd__nand2b_1 _08418_ (.A_N(\u_pwm.reg_ack_pwm2 ),
    .B(net1210),
    .Y(_03694_));
 sky130_fd_sc_hd__a22o_1 _08419_ (.A1(\u_pwm.reg_ack_pwm1 ),
    .A2(net1122),
    .B1(net1117),
    .B2(_03694_),
    .X(_03695_));
 sky130_fd_sc_hd__o21a_1 _08420_ (.A1(\u_pwm.reg_ack_pwm0 ),
    .A2(net1111),
    .B1(_03695_),
    .X(_03696_));
 sky130_fd_sc_hd__a21o_1 _08421_ (.A1(\u_pwm.reg_ack_glbl ),
    .A2(net1110),
    .B1(net1091),
    .X(_03697_));
 sky130_fd_sc_hd__o22a_1 _08422_ (.A1(\u_timer.reg_ack ),
    .A2(net723),
    .B1(_03696_),
    .B2(_03697_),
    .X(_03698_));
 sky130_fd_sc_hd__a22o_1 _08423_ (.A1(net1090),
    .A2(net65),
    .B1(net553),
    .B2(\u_ws281x.reg_ack ),
    .X(_03699_));
 sky130_fd_sc_hd__a221o_1 _08424_ (.A1(net2345),
    .A2(_03471_),
    .B1(_03698_),
    .B2(net559),
    .C1(_03699_),
    .X(_03700_));
 sky130_fd_sc_hd__and2_1 _08425_ (.A(\u_gpio.reg_ack ),
    .B(net548),
    .X(_03701_));
 sky130_fd_sc_hd__a211o_2 _08426_ (.A1(net1702),
    .A2(net544),
    .B1(net2346),
    .C1(_03701_),
    .X(net368));
 sky130_fd_sc_hd__o21a_1 _08427_ (.A1(net734),
    .A2(\u_ws281x.port0_rd ),
    .B1(_01195_),
    .X(_00621_));
 sky130_fd_sc_hd__a21oi_2 _08428_ (.A1(\u_ws281x.port0_enb ),
    .A2(_01177_),
    .B1(net2099),
    .Y(_03702_));
 sky130_fd_sc_hd__a31o_1 _08429_ (.A1(\u_ws281x.port0_enb ),
    .A2(_00825_),
    .A3(_01177_),
    .B1(_01196_),
    .X(_03703_));
 sky130_fd_sc_hd__and2_1 _08430_ (.A(_00798_),
    .B(net526),
    .X(_00605_));
 sky130_fd_sc_hd__o21ai_1 _08431_ (.A1(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .B1(net526),
    .Y(_03704_));
 sky130_fd_sc_hd__a21oi_1 _08432_ (.A1(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .B1(_03704_),
    .Y(_00612_));
 sky130_fd_sc_hd__and3_1 _08433_ (.A(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .C(\u_ws281x.u_txd_0.clk_cnt[2] ),
    .X(_03705_));
 sky130_fd_sc_hd__inv_2 _08434_ (.A(_03705_),
    .Y(_03706_));
 sky130_fd_sc_hd__a21o_1 _08435_ (.A1(\u_ws281x.u_txd_0.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_0.clk_cnt[1] ),
    .B1(\u_ws281x.u_txd_0.clk_cnt[2] ),
    .X(_03707_));
 sky130_fd_sc_hd__and3_1 _08436_ (.A(net526),
    .B(_03706_),
    .C(_03707_),
    .X(_00613_));
 sky130_fd_sc_hd__nor2_1 _08437_ (.A(_00804_),
    .B(_03706_),
    .Y(_03708_));
 sky130_fd_sc_hd__o21ai_1 _08438_ (.A1(\u_ws281x.u_txd_0.clk_cnt[3] ),
    .A2(_03705_),
    .B1(_03703_),
    .Y(_03709_));
 sky130_fd_sc_hd__nor2_1 _08439_ (.A(_03708_),
    .B(_03709_),
    .Y(_00614_));
 sky130_fd_sc_hd__and3_1 _08440_ (.A(\u_ws281x.u_txd_0.clk_cnt[3] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[4] ),
    .C(_03705_),
    .X(_03710_));
 sky130_fd_sc_hd__o21ai_1 _08441_ (.A1(\u_ws281x.u_txd_0.clk_cnt[4] ),
    .A2(_03708_),
    .B1(net526),
    .Y(_03711_));
 sky130_fd_sc_hd__nor2_1 _08442_ (.A(_03710_),
    .B(_03711_),
    .Y(_00615_));
 sky130_fd_sc_hd__and3_1 _08443_ (.A(\u_ws281x.u_txd_0.clk_cnt[4] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[5] ),
    .C(_03708_),
    .X(_03712_));
 sky130_fd_sc_hd__o21ai_1 _08444_ (.A1(\u_ws281x.u_txd_0.clk_cnt[5] ),
    .A2(_03710_),
    .B1(net526),
    .Y(_03713_));
 sky130_fd_sc_hd__nor2_1 _08445_ (.A(_03712_),
    .B(_03713_),
    .Y(_00616_));
 sky130_fd_sc_hd__and2_1 _08446_ (.A(\u_ws281x.u_txd_0.clk_cnt[6] ),
    .B(_03712_),
    .X(_03714_));
 sky130_fd_sc_hd__o21ai_1 _08447_ (.A1(\u_ws281x.u_txd_0.clk_cnt[6] ),
    .A2(_03712_),
    .B1(net526),
    .Y(_03715_));
 sky130_fd_sc_hd__nor2_1 _08448_ (.A(_03714_),
    .B(_03715_),
    .Y(_00617_));
 sky130_fd_sc_hd__and3_1 _08449_ (.A(\u_ws281x.u_txd_0.clk_cnt[6] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .C(_03712_),
    .X(_03716_));
 sky130_fd_sc_hd__o21ai_1 _08450_ (.A1(\u_ws281x.u_txd_0.clk_cnt[7] ),
    .A2(_03714_),
    .B1(net526),
    .Y(_03717_));
 sky130_fd_sc_hd__nor2_1 _08451_ (.A(_03716_),
    .B(_03717_),
    .Y(_00618_));
 sky130_fd_sc_hd__and2_1 _08452_ (.A(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .B(_03716_),
    .X(_03718_));
 sky130_fd_sc_hd__o21ai_1 _08453_ (.A1(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .A2(_03716_),
    .B1(net526),
    .Y(_03719_));
 sky130_fd_sc_hd__nor2_1 _08454_ (.A(_03718_),
    .B(_03719_),
    .Y(_00619_));
 sky130_fd_sc_hd__and3_1 _08455_ (.A(\u_ws281x.u_txd_0.clk_cnt[8] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .C(_03716_),
    .X(_03720_));
 sky130_fd_sc_hd__inv_2 _08456_ (.A(_03720_),
    .Y(_03721_));
 sky130_fd_sc_hd__o211a_1 _08457_ (.A1(\u_ws281x.u_txd_0.clk_cnt[9] ),
    .A2(_03718_),
    .B1(_03721_),
    .C1(net526),
    .X(_00620_));
 sky130_fd_sc_hd__nand2_1 _08458_ (.A(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .B(_03720_),
    .Y(_03722_));
 sky130_fd_sc_hd__o211a_1 _08459_ (.A1(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .A2(_03720_),
    .B1(_03722_),
    .C1(net526),
    .X(_00606_));
 sky130_fd_sc_hd__a21oi_1 _08460_ (.A1(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .A2(_03720_),
    .B1(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .Y(_03723_));
 sky130_fd_sc_hd__and3_1 _08461_ (.A(\u_ws281x.u_txd_0.clk_cnt[11] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[10] ),
    .C(_03720_),
    .X(_03724_));
 sky130_fd_sc_hd__nor3_1 _08462_ (.A(_03702_),
    .B(_03723_),
    .C(_03724_),
    .Y(_00607_));
 sky130_fd_sc_hd__and2_1 _08463_ (.A(\u_ws281x.u_txd_0.clk_cnt[12] ),
    .B(_03724_),
    .X(_03725_));
 sky130_fd_sc_hd__nor2_1 _08464_ (.A(\u_ws281x.u_txd_0.clk_cnt[12] ),
    .B(_03724_),
    .Y(_03726_));
 sky130_fd_sc_hd__nor3_1 _08465_ (.A(_03702_),
    .B(_03725_),
    .C(_03726_),
    .Y(_00608_));
 sky130_fd_sc_hd__a21oi_1 _08466_ (.A1(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .A2(_03725_),
    .B1(_03702_),
    .Y(_03727_));
 sky130_fd_sc_hd__o21a_1 _08467_ (.A1(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .A2(_03725_),
    .B1(_03727_),
    .X(_00609_));
 sky130_fd_sc_hd__a21oi_1 _08468_ (.A1(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .A2(_03725_),
    .B1(\u_ws281x.u_txd_0.clk_cnt[14] ),
    .Y(_03728_));
 sky130_fd_sc_hd__and3_1 _08469_ (.A(\u_ws281x.u_txd_0.clk_cnt[13] ),
    .B(\u_ws281x.u_txd_0.clk_cnt[14] ),
    .C(_03725_),
    .X(_03729_));
 sky130_fd_sc_hd__nor3_1 _08470_ (.A(_03702_),
    .B(_03728_),
    .C(_03729_),
    .Y(_00610_));
 sky130_fd_sc_hd__xnor2_1 _08471_ (.A(\u_ws281x.u_txd_0.clk_cnt[15] ),
    .B(_03729_),
    .Y(_03730_));
 sky130_fd_sc_hd__nor2_1 _08472_ (.A(_03702_),
    .B(_03730_),
    .Y(_00611_));
 sky130_fd_sc_hd__or2_1 _08473_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .B(_03376_),
    .X(_03731_));
 sky130_fd_sc_hd__o211a_1 _08474_ (.A1(net734),
    .A2(\u_ws281x.u_txd_0.led_data[0] ),
    .B1(net574),
    .C1(_03731_),
    .X(_00622_));
 sky130_fd_sc_hd__mux2_1 _08475_ (.A0(\u_ws281x.u_txd_0.led_data[1] ),
    .A1(_03381_),
    .S(net734),
    .X(_03732_));
 sky130_fd_sc_hd__mux2_1 _08476_ (.A0(\u_ws281x.u_txd_0.led_data[0] ),
    .A1(_03732_),
    .S(net574),
    .X(_00633_));
 sky130_fd_sc_hd__mux2_1 _08477_ (.A0(\u_ws281x.u_txd_0.led_data[2] ),
    .A1(_03387_),
    .S(net734),
    .X(_03733_));
 sky130_fd_sc_hd__mux2_1 _08478_ (.A0(\u_ws281x.u_txd_0.led_data[1] ),
    .A1(_03733_),
    .S(net574),
    .X(_00638_));
 sky130_fd_sc_hd__mux2_1 _08479_ (.A0(\u_ws281x.u_txd_0.led_data[3] ),
    .A1(_03391_),
    .S(net734),
    .X(_03734_));
 sky130_fd_sc_hd__mux2_1 _08480_ (.A0(\u_ws281x.u_txd_0.led_data[2] ),
    .A1(_03734_),
    .S(_01198_),
    .X(_00639_));
 sky130_fd_sc_hd__mux2_1 _08481_ (.A0(\u_ws281x.u_txd_0.led_data[4] ),
    .A1(_03395_),
    .S(net733),
    .X(_03735_));
 sky130_fd_sc_hd__mux2_1 _08482_ (.A0(\u_ws281x.u_txd_0.led_data[3] ),
    .A1(_03735_),
    .S(net573),
    .X(_00640_));
 sky130_fd_sc_hd__mux2_1 _08483_ (.A0(\u_ws281x.u_txd_0.led_data[5] ),
    .A1(_03399_),
    .S(net733),
    .X(_03736_));
 sky130_fd_sc_hd__mux2_1 _08484_ (.A0(\u_ws281x.u_txd_0.led_data[4] ),
    .A1(_03736_),
    .S(net573),
    .X(_00641_));
 sky130_fd_sc_hd__mux2_1 _08485_ (.A0(\u_ws281x.u_txd_0.led_data[6] ),
    .A1(_03403_),
    .S(net733),
    .X(_03737_));
 sky130_fd_sc_hd__mux2_1 _08486_ (.A0(\u_ws281x.u_txd_0.led_data[5] ),
    .A1(_03737_),
    .S(net573),
    .X(_00642_));
 sky130_fd_sc_hd__mux2_1 _08487_ (.A0(\u_ws281x.u_txd_0.led_data[7] ),
    .A1(_03406_),
    .S(net733),
    .X(_03738_));
 sky130_fd_sc_hd__mux2_1 _08488_ (.A0(\u_ws281x.u_txd_0.led_data[6] ),
    .A1(_03738_),
    .S(net573),
    .X(_00643_));
 sky130_fd_sc_hd__mux2_1 _08489_ (.A0(\u_ws281x.u_txd_0.led_data[8] ),
    .A1(_03408_),
    .S(net733),
    .X(_03739_));
 sky130_fd_sc_hd__mux2_1 _08490_ (.A0(\u_ws281x.u_txd_0.led_data[7] ),
    .A1(_03739_),
    .S(net573),
    .X(_00644_));
 sky130_fd_sc_hd__mux2_1 _08491_ (.A0(\u_ws281x.u_txd_0.led_data[9] ),
    .A1(_03411_),
    .S(net732),
    .X(_03740_));
 sky130_fd_sc_hd__mux2_1 _08492_ (.A0(\u_ws281x.u_txd_0.led_data[8] ),
    .A1(_03740_),
    .S(net571),
    .X(_00645_));
 sky130_fd_sc_hd__mux2_1 _08493_ (.A0(\u_ws281x.u_txd_0.led_data[10] ),
    .A1(_03414_),
    .S(net732),
    .X(_03741_));
 sky130_fd_sc_hd__mux2_1 _08494_ (.A0(\u_ws281x.u_txd_0.led_data[9] ),
    .A1(_03741_),
    .S(net571),
    .X(_00623_));
 sky130_fd_sc_hd__mux2_1 _08495_ (.A0(\u_ws281x.u_txd_0.led_data[11] ),
    .A1(_03418_),
    .S(net734),
    .X(_03742_));
 sky130_fd_sc_hd__mux2_1 _08496_ (.A0(\u_ws281x.u_txd_0.led_data[10] ),
    .A1(_03742_),
    .S(net572),
    .X(_00624_));
 sky130_fd_sc_hd__mux2_1 _08497_ (.A0(\u_ws281x.u_txd_0.led_data[12] ),
    .A1(_03421_),
    .S(net732),
    .X(_03743_));
 sky130_fd_sc_hd__mux2_1 _08498_ (.A0(\u_ws281x.u_txd_0.led_data[11] ),
    .A1(_03743_),
    .S(net572),
    .X(_00625_));
 sky130_fd_sc_hd__mux2_1 _08499_ (.A0(\u_ws281x.u_txd_0.led_data[13] ),
    .A1(_03424_),
    .S(net732),
    .X(_03744_));
 sky130_fd_sc_hd__mux2_1 _08500_ (.A0(\u_ws281x.u_txd_0.led_data[12] ),
    .A1(_03744_),
    .S(net572),
    .X(_00626_));
 sky130_fd_sc_hd__mux2_1 _08501_ (.A0(\u_ws281x.u_txd_0.led_data[14] ),
    .A1(_03426_),
    .S(net733),
    .X(_03745_));
 sky130_fd_sc_hd__mux2_1 _08502_ (.A0(\u_ws281x.u_txd_0.led_data[13] ),
    .A1(_03745_),
    .S(net572),
    .X(_00627_));
 sky130_fd_sc_hd__mux2_1 _08503_ (.A0(\u_ws281x.u_txd_0.led_data[15] ),
    .A1(_03429_),
    .S(net733),
    .X(_03746_));
 sky130_fd_sc_hd__mux2_1 _08504_ (.A0(\u_ws281x.u_txd_0.led_data[14] ),
    .A1(_03746_),
    .S(net571),
    .X(_00628_));
 sky130_fd_sc_hd__mux2_1 _08505_ (.A0(\u_ws281x.u_txd_0.led_data[16] ),
    .A1(_03433_),
    .S(net733),
    .X(_03747_));
 sky130_fd_sc_hd__mux2_1 _08506_ (.A0(\u_ws281x.u_txd_0.led_data[15] ),
    .A1(_03747_),
    .S(net571),
    .X(_00629_));
 sky130_fd_sc_hd__mux2_1 _08507_ (.A0(\u_ws281x.u_txd_0.led_data[17] ),
    .A1(_03436_),
    .S(net733),
    .X(_03748_));
 sky130_fd_sc_hd__mux2_1 _08508_ (.A0(\u_ws281x.u_txd_0.led_data[16] ),
    .A1(_03748_),
    .S(net571),
    .X(_00630_));
 sky130_fd_sc_hd__mux2_1 _08509_ (.A0(\u_ws281x.u_txd_0.led_data[18] ),
    .A1(_03438_),
    .S(net732),
    .X(_03749_));
 sky130_fd_sc_hd__mux2_1 _08510_ (.A0(\u_ws281x.u_txd_0.led_data[17] ),
    .A1(_03749_),
    .S(net571),
    .X(_00631_));
 sky130_fd_sc_hd__mux2_1 _08511_ (.A0(\u_ws281x.u_txd_0.led_data[19] ),
    .A1(_03442_),
    .S(net732),
    .X(_03750_));
 sky130_fd_sc_hd__mux2_1 _08512_ (.A0(\u_ws281x.u_txd_0.led_data[18] ),
    .A1(_03750_),
    .S(net571),
    .X(_00632_));
 sky130_fd_sc_hd__mux2_1 _08513_ (.A0(\u_ws281x.u_txd_0.led_data[20] ),
    .A1(_03444_),
    .S(net732),
    .X(_03751_));
 sky130_fd_sc_hd__mux2_1 _08514_ (.A0(\u_ws281x.u_txd_0.led_data[19] ),
    .A1(_03751_),
    .S(net571),
    .X(_00634_));
 sky130_fd_sc_hd__mux2_1 _08515_ (.A0(\u_ws281x.u_txd_0.led_data[21] ),
    .A1(_03448_),
    .S(net732),
    .X(_03752_));
 sky130_fd_sc_hd__mux2_1 _08516_ (.A0(\u_ws281x.u_txd_0.led_data[20] ),
    .A1(_03752_),
    .S(net571),
    .X(_00635_));
 sky130_fd_sc_hd__mux2_1 _08517_ (.A0(\u_ws281x.u_txd_0.led_data[22] ),
    .A1(_03450_),
    .S(net732),
    .X(_03753_));
 sky130_fd_sc_hd__mux2_1 _08518_ (.A0(\u_ws281x.u_txd_0.led_data[21] ),
    .A1(_03753_),
    .S(net571),
    .X(_00636_));
 sky130_fd_sc_hd__mux2_1 _08519_ (.A0(\u_ws281x.u_txd_0.led_data[23] ),
    .A1(_03454_),
    .S(net732),
    .X(_03754_));
 sky130_fd_sc_hd__mux2_1 _08520_ (.A0(\u_ws281x.u_txd_0.led_data[22] ),
    .A1(_03754_),
    .S(net572),
    .X(_00637_));
 sky130_fd_sc_hd__o21ai_1 _08521_ (.A1(net734),
    .A2(\u_ws281x.u_txd_0.bit_cnt[0] ),
    .B1(net574),
    .Y(_03755_));
 sky130_fd_sc_hd__o21ai_1 _08522_ (.A1(\u_ws281x.u_txd_0.bit_cnt[0] ),
    .A2(net574),
    .B1(_03755_),
    .Y(_00600_));
 sky130_fd_sc_hd__o21a_1 _08523_ (.A1(\u_ws281x.u_txd_0.bit_cnt[0] ),
    .A2(_00825_),
    .B1(\u_ws281x.u_txd_0.bit_cnt[1] ),
    .X(_03756_));
 sky130_fd_sc_hd__nor3_1 _08524_ (.A(\u_ws281x.u_txd_0.bit_cnt[0] ),
    .B(\u_ws281x.u_txd_0.bit_cnt[1] ),
    .C(net574),
    .Y(_03757_));
 sky130_fd_sc_hd__nor2_1 _08525_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .B(_01199_),
    .Y(_03758_));
 sky130_fd_sc_hd__or3_1 _08526_ (.A(_03756_),
    .B(_03757_),
    .C(_03758_),
    .X(_00601_));
 sky130_fd_sc_hd__nor3_1 _08527_ (.A(\u_ws281x.u_txd_0.bit_cnt[2] ),
    .B(_03757_),
    .C(_03758_),
    .Y(_03759_));
 sky130_fd_sc_hd__a21oi_1 _08528_ (.A1(\u_ws281x.u_txd_0.bit_cnt[2] ),
    .A2(_03757_),
    .B1(_03759_),
    .Y(_00602_));
 sky130_fd_sc_hd__xnor2_1 _08529_ (.A(\u_ws281x.u_txd_0.bit_cnt[3] ),
    .B(_01197_),
    .Y(_03760_));
 sky130_fd_sc_hd__a32o_1 _08530_ (.A1(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .A2(\u_ws281x.u_txd_0.bit_cnt[3] ),
    .A3(_00825_),
    .B1(_01199_),
    .B2(_03760_),
    .X(_00603_));
 sky130_fd_sc_hd__o31a_1 _08531_ (.A1(\u_ws281x.u_txd_0.bit_cnt[3] ),
    .A2(_00825_),
    .A3(_01197_),
    .B1(\u_ws281x.u_txd_0.bit_cnt[4] ),
    .X(_03761_));
 sky130_fd_sc_hd__or2_1 _08532_ (.A(_03758_),
    .B(_03761_),
    .X(_00604_));
 sky130_fd_sc_hd__o21a_1 _08533_ (.A1(net731),
    .A2(\u_ws281x.port1_rd ),
    .B1(_01237_),
    .X(_00672_));
 sky130_fd_sc_hd__o21a_1 _08534_ (.A1(_00838_),
    .A2(_01219_),
    .B1(_00839_),
    .X(_03762_));
 sky130_fd_sc_hd__o21ba_1 _08535_ (.A1(_00839_),
    .A2(_01236_),
    .B1_N(_03762_),
    .X(_03763_));
 sky130_fd_sc_hd__and2_1 _08536_ (.A(_00826_),
    .B(net525),
    .X(_00656_));
 sky130_fd_sc_hd__o21ai_1 _08537_ (.A1(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .B1(net525),
    .Y(_03764_));
 sky130_fd_sc_hd__a21oi_1 _08538_ (.A1(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .B1(_03764_),
    .Y(_00663_));
 sky130_fd_sc_hd__and3_1 _08539_ (.A(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .C(\u_ws281x.u_txd_1.clk_cnt[2] ),
    .X(_03765_));
 sky130_fd_sc_hd__inv_2 _08540_ (.A(_03765_),
    .Y(_03766_));
 sky130_fd_sc_hd__a21o_1 _08541_ (.A1(\u_ws281x.u_txd_1.clk_cnt[0] ),
    .A2(\u_ws281x.u_txd_1.clk_cnt[1] ),
    .B1(\u_ws281x.u_txd_1.clk_cnt[2] ),
    .X(_03767_));
 sky130_fd_sc_hd__and3_1 _08542_ (.A(net525),
    .B(_03766_),
    .C(_03767_),
    .X(_00664_));
 sky130_fd_sc_hd__nor2_1 _08543_ (.A(_00829_),
    .B(_03766_),
    .Y(_03768_));
 sky130_fd_sc_hd__o21ai_1 _08544_ (.A1(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .A2(_03765_),
    .B1(net525),
    .Y(_03769_));
 sky130_fd_sc_hd__nor2_1 _08545_ (.A(_03768_),
    .B(_03769_),
    .Y(_00665_));
 sky130_fd_sc_hd__and3_1 _08546_ (.A(\u_ws281x.u_txd_1.clk_cnt[3] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[4] ),
    .C(_03765_),
    .X(_03770_));
 sky130_fd_sc_hd__o21ai_1 _08547_ (.A1(\u_ws281x.u_txd_1.clk_cnt[4] ),
    .A2(_03768_),
    .B1(net525),
    .Y(_03771_));
 sky130_fd_sc_hd__nor2_1 _08548_ (.A(_03770_),
    .B(_03771_),
    .Y(_00666_));
 sky130_fd_sc_hd__and3_1 _08549_ (.A(\u_ws281x.u_txd_1.clk_cnt[4] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .C(_03768_),
    .X(_03772_));
 sky130_fd_sc_hd__o21ai_1 _08550_ (.A1(\u_ws281x.u_txd_1.clk_cnt[5] ),
    .A2(_03770_),
    .B1(_03763_),
    .Y(_03773_));
 sky130_fd_sc_hd__nor2_1 _08551_ (.A(_03772_),
    .B(_03773_),
    .Y(_00667_));
 sky130_fd_sc_hd__and2_1 _08552_ (.A(\u_ws281x.u_txd_1.clk_cnt[6] ),
    .B(_03772_),
    .X(_03774_));
 sky130_fd_sc_hd__o21ai_1 _08553_ (.A1(\u_ws281x.u_txd_1.clk_cnt[6] ),
    .A2(_03772_),
    .B1(net525),
    .Y(_03775_));
 sky130_fd_sc_hd__nor2_1 _08554_ (.A(_03774_),
    .B(_03775_),
    .Y(_00668_));
 sky130_fd_sc_hd__and3_1 _08555_ (.A(\u_ws281x.u_txd_1.clk_cnt[6] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .C(_03772_),
    .X(_03776_));
 sky130_fd_sc_hd__o21ai_1 _08556_ (.A1(\u_ws281x.u_txd_1.clk_cnt[7] ),
    .A2(_03774_),
    .B1(net525),
    .Y(_03777_));
 sky130_fd_sc_hd__nor2_1 _08557_ (.A(_03776_),
    .B(_03777_),
    .Y(_00669_));
 sky130_fd_sc_hd__and2_1 _08558_ (.A(\u_ws281x.u_txd_1.clk_cnt[8] ),
    .B(_03776_),
    .X(_03778_));
 sky130_fd_sc_hd__o21ai_1 _08559_ (.A1(\u_ws281x.u_txd_1.clk_cnt[8] ),
    .A2(_03776_),
    .B1(net525),
    .Y(_03779_));
 sky130_fd_sc_hd__nor2_1 _08560_ (.A(_03778_),
    .B(_03779_),
    .Y(_00670_));
 sky130_fd_sc_hd__and3_1 _08561_ (.A(\u_ws281x.u_txd_1.clk_cnt[8] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .C(_03776_),
    .X(_03780_));
 sky130_fd_sc_hd__inv_2 _08562_ (.A(_03780_),
    .Y(_03781_));
 sky130_fd_sc_hd__o211a_1 _08563_ (.A1(\u_ws281x.u_txd_1.clk_cnt[9] ),
    .A2(_03778_),
    .B1(_03781_),
    .C1(net525),
    .X(_00671_));
 sky130_fd_sc_hd__nand2_1 _08564_ (.A(\u_ws281x.u_txd_1.clk_cnt[10] ),
    .B(_03780_),
    .Y(_03782_));
 sky130_fd_sc_hd__o211a_1 _08565_ (.A1(\u_ws281x.u_txd_1.clk_cnt[10] ),
    .A2(_03780_),
    .B1(_03782_),
    .C1(net525),
    .X(_00657_));
 sky130_fd_sc_hd__nor2_1 _08566_ (.A(_00836_),
    .B(_03782_),
    .Y(_03783_));
 sky130_fd_sc_hd__or2_1 _08567_ (.A(_03762_),
    .B(_03783_),
    .X(_03784_));
 sky130_fd_sc_hd__a21oi_1 _08568_ (.A1(_00836_),
    .A2(_03782_),
    .B1(_03784_),
    .Y(_00658_));
 sky130_fd_sc_hd__and2_1 _08569_ (.A(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .B(_03783_),
    .X(_03785_));
 sky130_fd_sc_hd__nor2_1 _08570_ (.A(_03762_),
    .B(_03785_),
    .Y(_03786_));
 sky130_fd_sc_hd__o21a_1 _08571_ (.A1(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .A2(_03783_),
    .B1(_03786_),
    .X(_00659_));
 sky130_fd_sc_hd__and3_1 _08572_ (.A(\u_ws281x.u_txd_1.clk_cnt[13] ),
    .B(\u_ws281x.u_txd_1.clk_cnt[12] ),
    .C(_03783_),
    .X(_03787_));
 sky130_fd_sc_hd__nor2_1 _08573_ (.A(_03762_),
    .B(_03787_),
    .Y(_03788_));
 sky130_fd_sc_hd__o21a_1 _08574_ (.A1(\u_ws281x.u_txd_1.clk_cnt[13] ),
    .A2(_03785_),
    .B1(_03788_),
    .X(_00660_));
 sky130_fd_sc_hd__or2_1 _08575_ (.A(\u_ws281x.u_txd_1.clk_cnt[14] ),
    .B(_03787_),
    .X(_03789_));
 sky130_fd_sc_hd__nand2_1 _08576_ (.A(\u_ws281x.u_txd_1.clk_cnt[14] ),
    .B(_03787_),
    .Y(_03790_));
 sky130_fd_sc_hd__and3b_1 _08577_ (.A_N(_03762_),
    .B(_03789_),
    .C(_03790_),
    .X(_00661_));
 sky130_fd_sc_hd__or2_1 _08578_ (.A(\u_ws281x.u_txd_1.clk_cnt[15] ),
    .B(_03790_),
    .X(_03791_));
 sky130_fd_sc_hd__nand2_1 _08579_ (.A(\u_ws281x.u_txd_1.clk_cnt[15] ),
    .B(_03790_),
    .Y(_03792_));
 sky130_fd_sc_hd__a21oi_1 _08580_ (.A1(_03791_),
    .A2(_03792_),
    .B1(_03762_),
    .Y(_00662_));
 sky130_fd_sc_hd__or2_1 _08581_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .B(_03377_),
    .X(_03793_));
 sky130_fd_sc_hd__o211a_1 _08582_ (.A1(net731),
    .A2(\u_ws281x.u_txd_1.led_data[0] ),
    .B1(net570),
    .C1(_03793_),
    .X(_00673_));
 sky130_fd_sc_hd__mux2_1 _08583_ (.A0(\u_ws281x.u_txd_1.led_data[1] ),
    .A1(_03382_),
    .S(net731),
    .X(_03794_));
 sky130_fd_sc_hd__mux2_1 _08584_ (.A0(\u_ws281x.u_txd_1.led_data[0] ),
    .A1(_03794_),
    .S(net570),
    .X(_00684_));
 sky130_fd_sc_hd__mux2_1 _08585_ (.A0(\u_ws281x.u_txd_1.led_data[2] ),
    .A1(_03388_),
    .S(net731),
    .X(_03795_));
 sky130_fd_sc_hd__mux2_1 _08586_ (.A0(\u_ws281x.u_txd_1.led_data[1] ),
    .A1(_03795_),
    .S(net570),
    .X(_00689_));
 sky130_fd_sc_hd__mux2_1 _08587_ (.A0(\u_ws281x.u_txd_1.led_data[3] ),
    .A1(_03392_),
    .S(net731),
    .X(_03796_));
 sky130_fd_sc_hd__mux2_1 _08588_ (.A0(\u_ws281x.u_txd_1.led_data[2] ),
    .A1(_03796_),
    .S(net570),
    .X(_00690_));
 sky130_fd_sc_hd__mux2_1 _08589_ (.A0(\u_ws281x.u_txd_1.led_data[4] ),
    .A1(_03396_),
    .S(net731),
    .X(_03797_));
 sky130_fd_sc_hd__mux2_1 _08590_ (.A0(\u_ws281x.u_txd_1.led_data[3] ),
    .A1(_03797_),
    .S(net570),
    .X(_00691_));
 sky130_fd_sc_hd__mux2_1 _08591_ (.A0(\u_ws281x.u_txd_1.led_data[5] ),
    .A1(_03400_),
    .S(net731),
    .X(_03798_));
 sky130_fd_sc_hd__mux2_1 _08592_ (.A0(\u_ws281x.u_txd_1.led_data[4] ),
    .A1(_03798_),
    .S(net569),
    .X(_00692_));
 sky130_fd_sc_hd__mux2_1 _08593_ (.A0(\u_ws281x.u_txd_1.led_data[6] ),
    .A1(_03402_),
    .S(net731),
    .X(_03799_));
 sky130_fd_sc_hd__mux2_1 _08594_ (.A0(\u_ws281x.u_txd_1.led_data[5] ),
    .A1(_03799_),
    .S(net569),
    .X(_00693_));
 sky130_fd_sc_hd__mux2_1 _08595_ (.A0(\u_ws281x.u_txd_1.led_data[7] ),
    .A1(_03405_),
    .S(net731),
    .X(_03800_));
 sky130_fd_sc_hd__mux2_1 _08596_ (.A0(\u_ws281x.u_txd_1.led_data[6] ),
    .A1(_03800_),
    .S(net569),
    .X(_00694_));
 sky130_fd_sc_hd__mux2_1 _08597_ (.A0(\u_ws281x.u_txd_1.led_data[8] ),
    .A1(_03409_),
    .S(net730),
    .X(_03801_));
 sky130_fd_sc_hd__mux2_1 _08598_ (.A0(\u_ws281x.u_txd_1.led_data[7] ),
    .A1(_03801_),
    .S(net569),
    .X(_00695_));
 sky130_fd_sc_hd__mux2_1 _08599_ (.A0(\u_ws281x.u_txd_1.led_data[9] ),
    .A1(_03412_),
    .S(net730),
    .X(_03802_));
 sky130_fd_sc_hd__mux2_1 _08600_ (.A0(\u_ws281x.u_txd_1.led_data[8] ),
    .A1(_03802_),
    .S(net569),
    .X(_00696_));
 sky130_fd_sc_hd__mux2_1 _08601_ (.A0(\u_ws281x.u_txd_1.led_data[10] ),
    .A1(_03415_),
    .S(net730),
    .X(_03803_));
 sky130_fd_sc_hd__mux2_1 _08602_ (.A0(\u_ws281x.u_txd_1.led_data[9] ),
    .A1(_03803_),
    .S(net569),
    .X(_00674_));
 sky130_fd_sc_hd__mux2_1 _08603_ (.A0(\u_ws281x.u_txd_1.led_data[11] ),
    .A1(_03417_),
    .S(net730),
    .X(_03804_));
 sky130_fd_sc_hd__mux2_1 _08604_ (.A0(\u_ws281x.u_txd_1.led_data[10] ),
    .A1(_03804_),
    .S(net569),
    .X(_00675_));
 sky130_fd_sc_hd__mux2_1 _08605_ (.A0(\u_ws281x.u_txd_1.led_data[12] ),
    .A1(_03420_),
    .S(net730),
    .X(_03805_));
 sky130_fd_sc_hd__mux2_1 _08606_ (.A0(\u_ws281x.u_txd_1.led_data[11] ),
    .A1(_03805_),
    .S(net569),
    .X(_00676_));
 sky130_fd_sc_hd__mux2_1 _08607_ (.A0(\u_ws281x.u_txd_1.led_data[13] ),
    .A1(_03423_),
    .S(net729),
    .X(_03806_));
 sky130_fd_sc_hd__mux2_1 _08608_ (.A0(\u_ws281x.u_txd_1.led_data[12] ),
    .A1(_03806_),
    .S(net568),
    .X(_00677_));
 sky130_fd_sc_hd__mux2_1 _08609_ (.A0(\u_ws281x.u_txd_1.led_data[14] ),
    .A1(_03427_),
    .S(net729),
    .X(_03807_));
 sky130_fd_sc_hd__mux2_1 _08610_ (.A0(\u_ws281x.u_txd_1.led_data[13] ),
    .A1(_03807_),
    .S(net568),
    .X(_00678_));
 sky130_fd_sc_hd__mux2_1 _08611_ (.A0(\u_ws281x.u_txd_1.led_data[15] ),
    .A1(_03430_),
    .S(net730),
    .X(_03808_));
 sky130_fd_sc_hd__mux2_1 _08612_ (.A0(\u_ws281x.u_txd_1.led_data[14] ),
    .A1(_03808_),
    .S(net568),
    .X(_00679_));
 sky130_fd_sc_hd__mux2_1 _08613_ (.A0(\u_ws281x.u_txd_1.led_data[16] ),
    .A1(_03432_),
    .S(net729),
    .X(_03809_));
 sky130_fd_sc_hd__mux2_1 _08614_ (.A0(\u_ws281x.u_txd_1.led_data[15] ),
    .A1(_03809_),
    .S(net568),
    .X(_00680_));
 sky130_fd_sc_hd__mux2_1 _08615_ (.A0(\u_ws281x.u_txd_1.led_data[17] ),
    .A1(_03435_),
    .S(net729),
    .X(_03810_));
 sky130_fd_sc_hd__mux2_1 _08616_ (.A0(\u_ws281x.u_txd_1.led_data[16] ),
    .A1(_03810_),
    .S(net568),
    .X(_00681_));
 sky130_fd_sc_hd__mux2_1 _08617_ (.A0(\u_ws281x.u_txd_1.led_data[18] ),
    .A1(_03440_),
    .S(net729),
    .X(_03811_));
 sky130_fd_sc_hd__mux2_1 _08618_ (.A0(\u_ws281x.u_txd_1.led_data[17] ),
    .A1(_03811_),
    .S(net568),
    .X(_00682_));
 sky130_fd_sc_hd__mux2_1 _08619_ (.A0(\u_ws281x.u_txd_1.led_data[19] ),
    .A1(_03441_),
    .S(net729),
    .X(_03812_));
 sky130_fd_sc_hd__mux2_1 _08620_ (.A0(\u_ws281x.u_txd_1.led_data[18] ),
    .A1(_03812_),
    .S(net569),
    .X(_00683_));
 sky130_fd_sc_hd__mux2_1 _08621_ (.A0(\u_ws281x.u_txd_1.led_data[20] ),
    .A1(_03445_),
    .S(net729),
    .X(_03813_));
 sky130_fd_sc_hd__mux2_1 _08622_ (.A0(\u_ws281x.u_txd_1.led_data[19] ),
    .A1(_03813_),
    .S(net568),
    .X(_00685_));
 sky130_fd_sc_hd__mux2_1 _08623_ (.A0(\u_ws281x.u_txd_1.led_data[21] ),
    .A1(_03447_),
    .S(net729),
    .X(_03814_));
 sky130_fd_sc_hd__mux2_1 _08624_ (.A0(\u_ws281x.u_txd_1.led_data[20] ),
    .A1(_03814_),
    .S(net568),
    .X(_00686_));
 sky130_fd_sc_hd__mux2_1 _08625_ (.A0(\u_ws281x.u_txd_1.led_data[22] ),
    .A1(_03451_),
    .S(net729),
    .X(_03815_));
 sky130_fd_sc_hd__mux2_1 _08626_ (.A0(\u_ws281x.u_txd_1.led_data[21] ),
    .A1(_03815_),
    .S(net568),
    .X(_00687_));
 sky130_fd_sc_hd__mux2_1 _08627_ (.A0(\u_ws281x.u_txd_1.led_data[23] ),
    .A1(_03453_),
    .S(net729),
    .X(_03816_));
 sky130_fd_sc_hd__mux2_1 _08628_ (.A0(\u_ws281x.u_txd_1.led_data[22] ),
    .A1(_03816_),
    .S(net568),
    .X(_00688_));
 sky130_fd_sc_hd__o21ai_1 _08629_ (.A1(_00837_),
    .A2(\u_ws281x.u_txd_1.bit_cnt[0] ),
    .B1(_01239_),
    .Y(_03817_));
 sky130_fd_sc_hd__o21ai_1 _08630_ (.A1(\u_ws281x.u_txd_1.bit_cnt[0] ),
    .A2(net570),
    .B1(net2090),
    .Y(_00651_));
 sky130_fd_sc_hd__o21a_1 _08631_ (.A1(\u_ws281x.u_txd_1.bit_cnt[0] ),
    .A2(_00839_),
    .B1(\u_ws281x.u_txd_1.bit_cnt[1] ),
    .X(_03818_));
 sky130_fd_sc_hd__nor3_1 _08632_ (.A(\u_ws281x.u_txd_1.bit_cnt[0] ),
    .B(\u_ws281x.u_txd_1.bit_cnt[1] ),
    .C(net570),
    .Y(_03819_));
 sky130_fd_sc_hd__nor2_1 _08633_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .B(_01240_),
    .Y(_03820_));
 sky130_fd_sc_hd__or3_1 _08634_ (.A(_03818_),
    .B(_03819_),
    .C(_03820_),
    .X(_00652_));
 sky130_fd_sc_hd__nor3_1 _08635_ (.A(\u_ws281x.u_txd_1.bit_cnt[2] ),
    .B(_03819_),
    .C(_03820_),
    .Y(_03821_));
 sky130_fd_sc_hd__a21oi_1 _08636_ (.A1(\u_ws281x.u_txd_1.bit_cnt[2] ),
    .A2(_03819_),
    .B1(_03821_),
    .Y(_00653_));
 sky130_fd_sc_hd__xnor2_1 _08637_ (.A(\u_ws281x.u_txd_1.bit_cnt[3] ),
    .B(_01238_),
    .Y(_03822_));
 sky130_fd_sc_hd__a32o_1 _08638_ (.A1(net2247),
    .A2(\u_ws281x.u_txd_1.bit_cnt[3] ),
    .A3(_00839_),
    .B1(_01240_),
    .B2(_03822_),
    .X(_00654_));
 sky130_fd_sc_hd__o31a_1 _08639_ (.A1(\u_ws281x.u_txd_1.bit_cnt[3] ),
    .A2(_00839_),
    .A3(_01238_),
    .B1(\u_ws281x.u_txd_1.bit_cnt[4] ),
    .X(_03823_));
 sky130_fd_sc_hd__or2_1 _08640_ (.A(_03820_),
    .B(_03823_),
    .X(_00655_));
 sky130_fd_sc_hd__mux2_1 _08641_ (.A0(net2045),
    .A1(_00846_),
    .S(net522),
    .X(_00527_));
 sky130_fd_sc_hd__xnor2_1 _08642_ (.A(\u_timer.u_timer_0.timer_counter[0] ),
    .B(\u_timer.u_timer_0.timer_counter[1] ),
    .Y(_03824_));
 sky130_fd_sc_hd__mux2_1 _08643_ (.A0(net2064),
    .A1(_03824_),
    .S(net522),
    .X(_00534_));
 sky130_fd_sc_hd__o21ai_1 _08644_ (.A1(\u_timer.u_timer_0.timer_counter[0] ),
    .A2(\u_timer.u_timer_0.timer_counter[1] ),
    .B1(\u_timer.u_timer_0.timer_counter[2] ),
    .Y(_03825_));
 sky130_fd_sc_hd__nand2_1 _08645_ (.A(_01260_),
    .B(_03825_),
    .Y(_03826_));
 sky130_fd_sc_hd__mux2_1 _08646_ (.A0(net2061),
    .A1(_03826_),
    .S(net522),
    .X(_00535_));
 sky130_fd_sc_hd__nand2_1 _08647_ (.A(\u_timer.u_timer_0.timer_counter[3] ),
    .B(_01260_),
    .Y(_03827_));
 sky130_fd_sc_hd__nand2_1 _08648_ (.A(_01261_),
    .B(_03827_),
    .Y(_03828_));
 sky130_fd_sc_hd__mux2_1 _08649_ (.A0(net2053),
    .A1(_03828_),
    .S(net521),
    .X(_00536_));
 sky130_fd_sc_hd__xnor2_1 _08650_ (.A(\u_timer.u_timer_0.timer_counter[4] ),
    .B(_01261_),
    .Y(_03829_));
 sky130_fd_sc_hd__mux2_1 _08651_ (.A0(net2048),
    .A1(_03829_),
    .S(net522),
    .X(_00537_));
 sky130_fd_sc_hd__o21ai_1 _08652_ (.A1(\u_timer.u_timer_0.timer_counter[4] ),
    .A2(_01261_),
    .B1(\u_timer.u_timer_0.timer_counter[5] ),
    .Y(_03830_));
 sky130_fd_sc_hd__nand2_1 _08653_ (.A(_01262_),
    .B(_03830_),
    .Y(_03831_));
 sky130_fd_sc_hd__mux2_1 _08654_ (.A0(net2058),
    .A1(_03831_),
    .S(net522),
    .X(_00538_));
 sky130_fd_sc_hd__nand2_1 _08655_ (.A(\u_timer.u_timer_0.timer_counter[6] ),
    .B(_01262_),
    .Y(_03832_));
 sky130_fd_sc_hd__nand2_1 _08656_ (.A(_01263_),
    .B(_03832_),
    .Y(_03833_));
 sky130_fd_sc_hd__mux2_1 _08657_ (.A0(net2044),
    .A1(_03833_),
    .S(net522),
    .X(_00539_));
 sky130_fd_sc_hd__xnor2_1 _08658_ (.A(\u_timer.u_timer_0.timer_counter[7] ),
    .B(_01263_),
    .Y(_03834_));
 sky130_fd_sc_hd__mux2_1 _08659_ (.A0(net2042),
    .A1(_03834_),
    .S(net522),
    .X(_00540_));
 sky130_fd_sc_hd__o21ai_1 _08660_ (.A1(\u_timer.u_timer_0.timer_counter[7] ),
    .A2(_01263_),
    .B1(\u_timer.u_timer_0.timer_counter[8] ),
    .Y(_03835_));
 sky130_fd_sc_hd__nand2_1 _08661_ (.A(_01264_),
    .B(_03835_),
    .Y(_03836_));
 sky130_fd_sc_hd__mux2_1 _08662_ (.A0(net2324),
    .A1(_03836_),
    .S(net522),
    .X(_00541_));
 sky130_fd_sc_hd__nand2_1 _08663_ (.A(\u_timer.u_timer_0.timer_counter[9] ),
    .B(_01264_),
    .Y(_03837_));
 sky130_fd_sc_hd__nand2_1 _08664_ (.A(_01265_),
    .B(_03837_),
    .Y(_03838_));
 sky130_fd_sc_hd__mux2_1 _08665_ (.A0(net2328),
    .A1(_03838_),
    .S(net521),
    .X(_00542_));
 sky130_fd_sc_hd__xnor2_1 _08666_ (.A(\u_timer.u_timer_0.timer_counter[10] ),
    .B(_01265_),
    .Y(_03839_));
 sky130_fd_sc_hd__mux2_1 _08667_ (.A0(net2336),
    .A1(_03839_),
    .S(net521),
    .X(_00528_));
 sky130_fd_sc_hd__o21ai_1 _08668_ (.A1(\u_timer.u_timer_0.timer_counter[10] ),
    .A2(_01265_),
    .B1(\u_timer.u_timer_0.timer_counter[11] ),
    .Y(_03840_));
 sky130_fd_sc_hd__nand2_1 _08669_ (.A(_01266_),
    .B(_03840_),
    .Y(_03841_));
 sky130_fd_sc_hd__mux2_1 _08670_ (.A0(net2326),
    .A1(_03841_),
    .S(net521),
    .X(_00529_));
 sky130_fd_sc_hd__nand2_1 _08671_ (.A(\u_timer.u_timer_0.timer_counter[12] ),
    .B(_01266_),
    .Y(_03842_));
 sky130_fd_sc_hd__nand2_1 _08672_ (.A(_01267_),
    .B(_03842_),
    .Y(_03843_));
 sky130_fd_sc_hd__mux2_1 _08673_ (.A0(net2323),
    .A1(_03843_),
    .S(net521),
    .X(_00530_));
 sky130_fd_sc_hd__xnor2_1 _08674_ (.A(\u_timer.u_timer_0.timer_counter[13] ),
    .B(_01267_),
    .Y(_03844_));
 sky130_fd_sc_hd__mux2_1 _08675_ (.A0(net2332),
    .A1(_03844_),
    .S(net521),
    .X(_00531_));
 sky130_fd_sc_hd__o21ai_1 _08676_ (.A1(\u_timer.u_timer_0.timer_counter[13] ),
    .A2(_01267_),
    .B1(\u_timer.u_timer_0.timer_counter[14] ),
    .Y(_03845_));
 sky130_fd_sc_hd__nand2_1 _08677_ (.A(_01268_),
    .B(_03845_),
    .Y(_03846_));
 sky130_fd_sc_hd__mux2_1 _08678_ (.A0(net2310),
    .A1(_03846_),
    .S(net521),
    .X(_00532_));
 sky130_fd_sc_hd__and2_1 _08679_ (.A(\u_timer.u_timer_0.timer_counter[15] ),
    .B(_01268_),
    .X(_03847_));
 sky130_fd_sc_hd__or3b_1 _08680_ (.A(\u_timer.u_timer_0.timer_hit ),
    .B(_03847_),
    .C_N(net521),
    .X(_03848_));
 sky130_fd_sc_hd__o21a_1 _08681_ (.A1(net2337),
    .A2(net521),
    .B1(_03848_),
    .X(_00533_));
 sky130_fd_sc_hd__mux2_1 _08682_ (.A0(net2330),
    .A1(_00843_),
    .S(net520),
    .X(_00544_));
 sky130_fd_sc_hd__xnor2_1 _08683_ (.A(\u_timer.u_timer_1.timer_counter[0] ),
    .B(\u_timer.u_timer_1.timer_counter[1] ),
    .Y(_03849_));
 sky130_fd_sc_hd__mux2_1 _08684_ (.A0(net2309),
    .A1(_03849_),
    .S(net520),
    .X(_00551_));
 sky130_fd_sc_hd__o21ai_1 _08685_ (.A1(\u_timer.u_timer_1.timer_counter[0] ),
    .A2(\u_timer.u_timer_1.timer_counter[1] ),
    .B1(\u_timer.u_timer_1.timer_counter[2] ),
    .Y(_03850_));
 sky130_fd_sc_hd__nand2_1 _08686_ (.A(_01251_),
    .B(_03850_),
    .Y(_03851_));
 sky130_fd_sc_hd__mux2_1 _08687_ (.A0(net2322),
    .A1(_03851_),
    .S(net520),
    .X(_00552_));
 sky130_fd_sc_hd__nand2_1 _08688_ (.A(\u_timer.u_timer_1.timer_counter[3] ),
    .B(_01251_),
    .Y(_03852_));
 sky130_fd_sc_hd__nand2_1 _08689_ (.A(_01252_),
    .B(_03852_),
    .Y(_03853_));
 sky130_fd_sc_hd__mux2_1 _08690_ (.A0(net2253),
    .A1(_03853_),
    .S(net520),
    .X(_00553_));
 sky130_fd_sc_hd__xnor2_1 _08691_ (.A(\u_timer.u_timer_1.timer_counter[4] ),
    .B(_01252_),
    .Y(_03854_));
 sky130_fd_sc_hd__mux2_1 _08692_ (.A0(net2242),
    .A1(_03854_),
    .S(net520),
    .X(_00554_));
 sky130_fd_sc_hd__o21ai_1 _08693_ (.A1(\u_timer.u_timer_1.timer_counter[4] ),
    .A2(_01252_),
    .B1(\u_timer.u_timer_1.timer_counter[5] ),
    .Y(_03855_));
 sky130_fd_sc_hd__nand2_1 _08694_ (.A(_01253_),
    .B(_03855_),
    .Y(_03856_));
 sky130_fd_sc_hd__mux2_1 _08695_ (.A0(net2244),
    .A1(_03856_),
    .S(net520),
    .X(_00555_));
 sky130_fd_sc_hd__nand2_1 _08696_ (.A(\u_timer.u_timer_1.timer_counter[6] ),
    .B(_01253_),
    .Y(_03857_));
 sky130_fd_sc_hd__nand2_1 _08697_ (.A(_01254_),
    .B(_03857_),
    .Y(_03858_));
 sky130_fd_sc_hd__mux2_1 _08698_ (.A0(net2261),
    .A1(_03858_),
    .S(net520),
    .X(_00556_));
 sky130_fd_sc_hd__xnor2_1 _08699_ (.A(\u_timer.u_timer_1.timer_counter[7] ),
    .B(_01254_),
    .Y(_03859_));
 sky130_fd_sc_hd__mux2_1 _08700_ (.A0(net2239),
    .A1(_03859_),
    .S(net520),
    .X(_00557_));
 sky130_fd_sc_hd__o21ai_1 _08701_ (.A1(\u_timer.u_timer_1.timer_counter[7] ),
    .A2(_01254_),
    .B1(\u_timer.u_timer_1.timer_counter[8] ),
    .Y(_03860_));
 sky130_fd_sc_hd__nand2_1 _08702_ (.A(_01255_),
    .B(_03860_),
    .Y(_03861_));
 sky130_fd_sc_hd__mux2_1 _08703_ (.A0(net2022),
    .A1(_03861_),
    .S(net519),
    .X(_00558_));
 sky130_fd_sc_hd__nand2_1 _08704_ (.A(\u_timer.u_timer_1.timer_counter[9] ),
    .B(_01255_),
    .Y(_03862_));
 sky130_fd_sc_hd__nand2_1 _08705_ (.A(_01256_),
    .B(_03862_),
    .Y(_03863_));
 sky130_fd_sc_hd__mux2_1 _08706_ (.A0(net2021),
    .A1(_03863_),
    .S(net519),
    .X(_00559_));
 sky130_fd_sc_hd__xnor2_1 _08707_ (.A(\u_timer.u_timer_1.timer_counter[10] ),
    .B(_01256_),
    .Y(_03864_));
 sky130_fd_sc_hd__mux2_1 _08708_ (.A0(net2023),
    .A1(_03864_),
    .S(net519),
    .X(_00545_));
 sky130_fd_sc_hd__o21ai_1 _08709_ (.A1(\u_timer.u_timer_1.timer_counter[10] ),
    .A2(_01256_),
    .B1(\u_timer.u_timer_1.timer_counter[11] ),
    .Y(_03865_));
 sky130_fd_sc_hd__nand2_1 _08710_ (.A(_01257_),
    .B(_03865_),
    .Y(_03866_));
 sky130_fd_sc_hd__mux2_1 _08711_ (.A0(net2024),
    .A1(_03866_),
    .S(net519),
    .X(_00546_));
 sky130_fd_sc_hd__nand2_1 _08712_ (.A(\u_timer.u_timer_1.timer_counter[12] ),
    .B(_01257_),
    .Y(_03867_));
 sky130_fd_sc_hd__nand2_1 _08713_ (.A(_01258_),
    .B(_03867_),
    .Y(_03868_));
 sky130_fd_sc_hd__mux2_1 _08714_ (.A0(net2039),
    .A1(_03868_),
    .S(net519),
    .X(_00547_));
 sky130_fd_sc_hd__xnor2_1 _08715_ (.A(\u_timer.u_timer_1.timer_counter[13] ),
    .B(_01258_),
    .Y(_03869_));
 sky130_fd_sc_hd__mux2_1 _08716_ (.A0(net2034),
    .A1(_03869_),
    .S(net519),
    .X(_00548_));
 sky130_fd_sc_hd__o21ai_1 _08717_ (.A1(\u_timer.u_timer_1.timer_counter[13] ),
    .A2(_01258_),
    .B1(\u_timer.u_timer_1.timer_counter[14] ),
    .Y(_03870_));
 sky130_fd_sc_hd__nand2_1 _08718_ (.A(_01259_),
    .B(_03870_),
    .Y(_03871_));
 sky130_fd_sc_hd__mux2_1 _08719_ (.A0(net2017),
    .A1(_03871_),
    .S(net519),
    .X(_00549_));
 sky130_fd_sc_hd__and2_1 _08720_ (.A(\u_timer.u_timer_1.timer_counter[15] ),
    .B(_01259_),
    .X(_03872_));
 sky130_fd_sc_hd__or3b_1 _08721_ (.A(\u_timer.u_timer_1.timer_hit ),
    .B(_03872_),
    .C_N(net519),
    .X(_03873_));
 sky130_fd_sc_hd__o21a_1 _08722_ (.A1(net2038),
    .A2(net519),
    .B1(_03873_),
    .X(_00550_));
 sky130_fd_sc_hd__mux2_1 _08723_ (.A0(net2250),
    .A1(_00840_),
    .S(net516),
    .X(_00561_));
 sky130_fd_sc_hd__xnor2_1 _08724_ (.A(\u_timer.u_timer_2.timer_counter[0] ),
    .B(\u_timer.u_timer_2.timer_counter[1] ),
    .Y(_03874_));
 sky130_fd_sc_hd__mux2_1 _08725_ (.A0(net2228),
    .A1(_03874_),
    .S(net516),
    .X(_00568_));
 sky130_fd_sc_hd__o21ai_1 _08726_ (.A1(\u_timer.u_timer_2.timer_counter[0] ),
    .A2(\u_timer.u_timer_2.timer_counter[1] ),
    .B1(\u_timer.u_timer_2.timer_counter[2] ),
    .Y(_03875_));
 sky130_fd_sc_hd__nand2_1 _08727_ (.A(_01242_),
    .B(_03875_),
    .Y(_03876_));
 sky130_fd_sc_hd__mux2_1 _08728_ (.A0(net2258),
    .A1(_03876_),
    .S(net516),
    .X(_00569_));
 sky130_fd_sc_hd__nand2_1 _08729_ (.A(\u_timer.u_timer_2.timer_counter[3] ),
    .B(_01242_),
    .Y(_03877_));
 sky130_fd_sc_hd__nand2_1 _08730_ (.A(_01243_),
    .B(_03877_),
    .Y(_03878_));
 sky130_fd_sc_hd__mux2_1 _08731_ (.A0(net2307),
    .A1(_03878_),
    .S(net516),
    .X(_00570_));
 sky130_fd_sc_hd__xnor2_1 _08732_ (.A(\u_timer.u_timer_2.timer_counter[4] ),
    .B(_01243_),
    .Y(_03879_));
 sky130_fd_sc_hd__mux2_1 _08733_ (.A0(net2269),
    .A1(_03879_),
    .S(net516),
    .X(_00571_));
 sky130_fd_sc_hd__o21ai_1 _08734_ (.A1(\u_timer.u_timer_2.timer_counter[4] ),
    .A2(_01243_),
    .B1(\u_timer.u_timer_2.timer_counter[5] ),
    .Y(_03880_));
 sky130_fd_sc_hd__nand2_1 _08735_ (.A(_01244_),
    .B(_03880_),
    .Y(_03881_));
 sky130_fd_sc_hd__mux2_1 _08736_ (.A0(net2251),
    .A1(_03881_),
    .S(net516),
    .X(_00572_));
 sky130_fd_sc_hd__nand2_1 _08737_ (.A(\u_timer.u_timer_2.timer_counter[6] ),
    .B(_01244_),
    .Y(_03882_));
 sky130_fd_sc_hd__nand2_1 _08738_ (.A(_01245_),
    .B(_03882_),
    .Y(_03883_));
 sky130_fd_sc_hd__mux2_1 _08739_ (.A0(net2263),
    .A1(_03883_),
    .S(net516),
    .X(_00573_));
 sky130_fd_sc_hd__xnor2_1 _08740_ (.A(\u_timer.u_timer_2.timer_counter[7] ),
    .B(_01245_),
    .Y(_03884_));
 sky130_fd_sc_hd__mux2_1 _08741_ (.A0(net2270),
    .A1(_03884_),
    .S(net515),
    .X(_00574_));
 sky130_fd_sc_hd__o21ai_1 _08742_ (.A1(\u_timer.u_timer_2.timer_counter[7] ),
    .A2(_01245_),
    .B1(\u_timer.u_timer_2.timer_counter[8] ),
    .Y(_03885_));
 sky130_fd_sc_hd__nand2_1 _08743_ (.A(_01246_),
    .B(_03885_),
    .Y(_03886_));
 sky130_fd_sc_hd__mux2_1 _08744_ (.A0(net2290),
    .A1(_03886_),
    .S(net515),
    .X(_00575_));
 sky130_fd_sc_hd__nand2_1 _08745_ (.A(\u_timer.u_timer_2.timer_counter[9] ),
    .B(_01246_),
    .Y(_03887_));
 sky130_fd_sc_hd__nand2_1 _08746_ (.A(_01247_),
    .B(_03887_),
    .Y(_03888_));
 sky130_fd_sc_hd__mux2_1 _08747_ (.A0(net2291),
    .A1(_03888_),
    .S(net516),
    .X(_00576_));
 sky130_fd_sc_hd__xnor2_1 _08748_ (.A(\u_timer.u_timer_2.timer_counter[10] ),
    .B(_01247_),
    .Y(_03889_));
 sky130_fd_sc_hd__mux2_1 _08749_ (.A0(net2298),
    .A1(_03889_),
    .S(net515),
    .X(_00562_));
 sky130_fd_sc_hd__o21ai_1 _08750_ (.A1(\u_timer.u_timer_2.timer_counter[10] ),
    .A2(_01247_),
    .B1(\u_timer.u_timer_2.timer_counter[11] ),
    .Y(_03890_));
 sky130_fd_sc_hd__nand2_1 _08751_ (.A(_01248_),
    .B(_03890_),
    .Y(_03891_));
 sky130_fd_sc_hd__mux2_1 _08752_ (.A0(net2308),
    .A1(_03891_),
    .S(net515),
    .X(_00563_));
 sky130_fd_sc_hd__nand2_1 _08753_ (.A(\u_timer.u_timer_2.timer_counter[12] ),
    .B(_01248_),
    .Y(_03892_));
 sky130_fd_sc_hd__nand2_1 _08754_ (.A(_01249_),
    .B(_03892_),
    .Y(_03893_));
 sky130_fd_sc_hd__mux2_1 _08755_ (.A0(net2288),
    .A1(_03893_),
    .S(net515),
    .X(_00564_));
 sky130_fd_sc_hd__xnor2_1 _08756_ (.A(\u_timer.u_timer_2.timer_counter[13] ),
    .B(_01249_),
    .Y(_03894_));
 sky130_fd_sc_hd__mux2_1 _08757_ (.A0(net2280),
    .A1(_03894_),
    .S(net515),
    .X(_00565_));
 sky130_fd_sc_hd__o21ai_1 _08758_ (.A1(\u_timer.u_timer_2.timer_counter[13] ),
    .A2(_01249_),
    .B1(\u_timer.u_timer_2.timer_counter[14] ),
    .Y(_03895_));
 sky130_fd_sc_hd__nand2_1 _08759_ (.A(_01250_),
    .B(_03895_),
    .Y(_03896_));
 sky130_fd_sc_hd__mux2_1 _08760_ (.A0(net2316),
    .A1(_03896_),
    .S(net515),
    .X(_00566_));
 sky130_fd_sc_hd__and2_1 _08761_ (.A(\u_timer.u_timer_2.timer_counter[15] ),
    .B(_01250_),
    .X(_03897_));
 sky130_fd_sc_hd__or3b_1 _08762_ (.A(\u_timer.u_timer_2.timer_hit ),
    .B(_03897_),
    .C_N(net515),
    .X(_03898_));
 sky130_fd_sc_hd__o21a_1 _08763_ (.A1(net2311),
    .A2(net515),
    .B1(_03898_),
    .X(_00567_));
 sky130_fd_sc_hd__and3_1 _08764_ (.A(\u_timer.u_pulse_1ms.cnt[1] ),
    .B(\u_timer.u_pulse_1ms.cnt[0] ),
    .C(\u_timer.u_pulse_1ms.cnt[2] ),
    .X(_03899_));
 sky130_fd_sc_hd__or2_1 _08765_ (.A(\u_timer.u_pulse_1ms.cnt[3] ),
    .B(_03899_),
    .X(_03900_));
 sky130_fd_sc_hd__and4_1 _08766_ (.A(\u_timer.u_pulse_1ms.cnt[5] ),
    .B(\u_timer.u_pulse_1ms.cnt[7] ),
    .C(\u_timer.u_pulse_1ms.cnt[6] ),
    .D(\u_timer.u_pulse_1ms.cnt[8] ),
    .X(_03901_));
 sky130_fd_sc_hd__o211ai_4 _08767_ (.A1(\u_timer.u_pulse_1ms.cnt[4] ),
    .A2(_03900_),
    .B1(_03901_),
    .C1(\u_timer.u_pulse_1ms.cnt[9] ),
    .Y(_03902_));
 sky130_fd_sc_hd__and2b_1 _08768_ (.A_N(\u_timer.u_pulse_1ms.cnt[0] ),
    .B(_03902_),
    .X(_00479_));
 sky130_fd_sc_hd__o21ai_1 _08769_ (.A1(\u_timer.u_pulse_1ms.cnt[1] ),
    .A2(\u_timer.u_pulse_1ms.cnt[0] ),
    .B1(_03902_),
    .Y(_03903_));
 sky130_fd_sc_hd__a21oi_1 _08770_ (.A1(\u_timer.u_pulse_1ms.cnt[1] ),
    .A2(\u_timer.u_pulse_1ms.cnt[0] ),
    .B1(_03903_),
    .Y(_00480_));
 sky130_fd_sc_hd__a21o_1 _08771_ (.A1(\u_timer.u_pulse_1ms.cnt[1] ),
    .A2(\u_timer.u_pulse_1ms.cnt[0] ),
    .B1(\u_timer.u_pulse_1ms.cnt[2] ),
    .X(_03904_));
 sky130_fd_sc_hd__and3b_1 _08772_ (.A_N(_03899_),
    .B(_03902_),
    .C(_03904_),
    .X(_00481_));
 sky130_fd_sc_hd__nand2_1 _08773_ (.A(\u_timer.u_pulse_1ms.cnt[3] ),
    .B(_03899_),
    .Y(_03905_));
 sky130_fd_sc_hd__and3_1 _08774_ (.A(_03900_),
    .B(_03902_),
    .C(_03905_),
    .X(_00482_));
 sky130_fd_sc_hd__a21o_1 _08775_ (.A1(\u_timer.u_pulse_1ms.cnt[3] ),
    .A2(_03899_),
    .B1(\u_timer.u_pulse_1ms.cnt[4] ),
    .X(_03906_));
 sky130_fd_sc_hd__and3_1 _08776_ (.A(\u_timer.u_pulse_1ms.cnt[3] ),
    .B(\u_timer.u_pulse_1ms.cnt[4] ),
    .C(_03899_),
    .X(_03907_));
 sky130_fd_sc_hd__clkinv_2 _08777_ (.A(_03907_),
    .Y(_03908_));
 sky130_fd_sc_hd__and3_1 _08778_ (.A(_03902_),
    .B(_03906_),
    .C(_03908_),
    .X(_00483_));
 sky130_fd_sc_hd__and2_1 _08779_ (.A(\u_timer.u_pulse_1ms.cnt[5] ),
    .B(_03907_),
    .X(_03909_));
 sky130_fd_sc_hd__o21ai_1 _08780_ (.A1(\u_timer.u_pulse_1ms.cnt[5] ),
    .A2(_03907_),
    .B1(_03902_),
    .Y(_03910_));
 sky130_fd_sc_hd__nor2_1 _08781_ (.A(_03909_),
    .B(_03910_),
    .Y(_00484_));
 sky130_fd_sc_hd__and3_1 _08782_ (.A(\u_timer.u_pulse_1ms.cnt[5] ),
    .B(\u_timer.u_pulse_1ms.cnt[6] ),
    .C(_03907_),
    .X(_03911_));
 sky130_fd_sc_hd__o21ai_1 _08783_ (.A1(\u_timer.u_pulse_1ms.cnt[6] ),
    .A2(_03909_),
    .B1(_03902_),
    .Y(_03912_));
 sky130_fd_sc_hd__nor2_1 _08784_ (.A(_03911_),
    .B(_03912_),
    .Y(_00485_));
 sky130_fd_sc_hd__and2_1 _08785_ (.A(\u_timer.u_pulse_1ms.cnt[7] ),
    .B(_03911_),
    .X(_03913_));
 sky130_fd_sc_hd__o21ai_1 _08786_ (.A1(\u_timer.u_pulse_1ms.cnt[7] ),
    .A2(_03911_),
    .B1(_03902_),
    .Y(_03914_));
 sky130_fd_sc_hd__nor2_1 _08787_ (.A(_03913_),
    .B(_03914_),
    .Y(_00486_));
 sky130_fd_sc_hd__nand2_1 _08788_ (.A(\u_timer.u_pulse_1ms.cnt[8] ),
    .B(_03913_),
    .Y(_03915_));
 sky130_fd_sc_hd__o211a_1 _08789_ (.A1(\u_timer.u_pulse_1ms.cnt[8] ),
    .A2(_03913_),
    .B1(_03915_),
    .C1(_03902_),
    .X(_00487_));
 sky130_fd_sc_hd__a21boi_1 _08790_ (.A1(_00856_),
    .A2(_03915_),
    .B1_N(_03902_),
    .Y(_00488_));
 sky130_fd_sc_hd__and3_1 _08791_ (.A(\u_timer.u_pulse_1s.cnt[7] ),
    .B(\u_timer.u_pulse_1s.cnt[6] ),
    .C(\u_timer.u_pulse_1s.cnt[8] ),
    .X(_03916_));
 sky130_fd_sc_hd__and3_1 _08792_ (.A(\u_timer.u_pulse_1s.cnt[5] ),
    .B(\u_timer.u_pulse_1s.cnt[9] ),
    .C(_03916_),
    .X(_03917_));
 sky130_fd_sc_hd__nand2_1 _08793_ (.A(\u_timer.u_pulse_1s.cnt[1] ),
    .B(\u_timer.u_pulse_1s.cnt[0] ),
    .Y(_03918_));
 sky130_fd_sc_hd__and3_2 _08794_ (.A(\u_timer.u_pulse_1s.cnt[1] ),
    .B(\u_timer.u_pulse_1s.cnt[0] ),
    .C(\u_timer.u_pulse_1s.cnt[2] ),
    .X(_03919_));
 sky130_fd_sc_hd__o31ai_4 _08795_ (.A1(\u_timer.u_pulse_1s.cnt[3] ),
    .A2(\u_timer.u_pulse_1s.cnt[4] ),
    .A3(_03919_),
    .B1(_03917_),
    .Y(_03920_));
 sky130_fd_sc_hd__and2b_1 _08796_ (.A_N(\u_timer.u_pulse_1s.cnt[0] ),
    .B(_03920_),
    .X(_00489_));
 sky130_fd_sc_hd__and3_1 _08797_ (.A(_01338_),
    .B(_03918_),
    .C(_03920_),
    .X(_00490_));
 sky130_fd_sc_hd__a21o_1 _08798_ (.A1(\u_timer.u_pulse_1s.cnt[1] ),
    .A2(\u_timer.u_pulse_1s.cnt[0] ),
    .B1(\u_timer.u_pulse_1s.cnt[2] ),
    .X(_03921_));
 sky130_fd_sc_hd__and3b_1 _08799_ (.A_N(_03919_),
    .B(_03920_),
    .C(_03921_),
    .X(_00491_));
 sky130_fd_sc_hd__a21oi_1 _08800_ (.A1(\u_timer.u_pulse_1s.cnt[3] ),
    .A2(_03919_),
    .B1(_03917_),
    .Y(_03922_));
 sky130_fd_sc_hd__o21a_1 _08801_ (.A1(\u_timer.u_pulse_1s.cnt[3] ),
    .A2(_03919_),
    .B1(_03922_),
    .X(_00492_));
 sky130_fd_sc_hd__a21oi_1 _08802_ (.A1(\u_timer.u_pulse_1s.cnt[3] ),
    .A2(_03919_),
    .B1(\u_timer.u_pulse_1s.cnt[4] ),
    .Y(_03923_));
 sky130_fd_sc_hd__and3_1 _08803_ (.A(\u_timer.u_pulse_1s.cnt[3] ),
    .B(\u_timer.u_pulse_1s.cnt[4] ),
    .C(_03919_),
    .X(_03924_));
 sky130_fd_sc_hd__nor3_1 _08804_ (.A(_03917_),
    .B(_03923_),
    .C(_03924_),
    .Y(_00493_));
 sky130_fd_sc_hd__and2_1 _08805_ (.A(\u_timer.u_pulse_1s.cnt[5] ),
    .B(_03924_),
    .X(_03925_));
 sky130_fd_sc_hd__o21ai_1 _08806_ (.A1(\u_timer.u_pulse_1s.cnt[5] ),
    .A2(_03924_),
    .B1(_03920_),
    .Y(_03926_));
 sky130_fd_sc_hd__nor2_1 _08807_ (.A(_03925_),
    .B(_03926_),
    .Y(_00494_));
 sky130_fd_sc_hd__and3_1 _08808_ (.A(\u_timer.u_pulse_1s.cnt[5] ),
    .B(\u_timer.u_pulse_1s.cnt[6] ),
    .C(_03924_),
    .X(_03927_));
 sky130_fd_sc_hd__o21ai_1 _08809_ (.A1(\u_timer.u_pulse_1s.cnt[6] ),
    .A2(_03925_),
    .B1(_03920_),
    .Y(_03928_));
 sky130_fd_sc_hd__nor2_1 _08810_ (.A(_03927_),
    .B(_03928_),
    .Y(_00495_));
 sky130_fd_sc_hd__and2_1 _08811_ (.A(\u_timer.u_pulse_1s.cnt[7] ),
    .B(_03927_),
    .X(_03929_));
 sky130_fd_sc_hd__o21ai_1 _08812_ (.A1(\u_timer.u_pulse_1s.cnt[7] ),
    .A2(_03927_),
    .B1(_03920_),
    .Y(_03930_));
 sky130_fd_sc_hd__nor2_1 _08813_ (.A(_03929_),
    .B(_03930_),
    .Y(_00496_));
 sky130_fd_sc_hd__nand2_1 _08814_ (.A(\u_timer.u_pulse_1s.cnt[8] ),
    .B(_03929_),
    .Y(_03931_));
 sky130_fd_sc_hd__o211a_1 _08815_ (.A1(\u_timer.u_pulse_1s.cnt[8] ),
    .A2(_03929_),
    .B1(_03931_),
    .C1(_03920_),
    .X(_00497_));
 sky130_fd_sc_hd__a21boi_1 _08816_ (.A1(_00857_),
    .A2(_03931_),
    .B1_N(_03920_),
    .Y(_00498_));
 sky130_fd_sc_hd__nor2_1 _08817_ (.A(\u_timer.u_pulse_1us.cnt[0] ),
    .B(_00499_),
    .Y(_00500_));
 sky130_fd_sc_hd__o21ai_1 _08818_ (.A1(\u_timer.u_pulse_1us.cnt[0] ),
    .A2(\u_timer.u_pulse_1us.cnt[1] ),
    .B1(_01531_),
    .Y(_03932_));
 sky130_fd_sc_hd__a21oi_1 _08819_ (.A1(\u_timer.u_pulse_1us.cnt[0] ),
    .A2(\u_timer.u_pulse_1us.cnt[1] ),
    .B1(_03932_),
    .Y(_00501_));
 sky130_fd_sc_hd__and3_1 _08820_ (.A(\u_timer.u_pulse_1us.cnt[0] ),
    .B(\u_timer.u_pulse_1us.cnt[1] ),
    .C(\u_timer.u_pulse_1us.cnt[2] ),
    .X(_03933_));
 sky130_fd_sc_hd__inv_2 _08821_ (.A(_03933_),
    .Y(_03934_));
 sky130_fd_sc_hd__a21o_1 _08822_ (.A1(\u_timer.u_pulse_1us.cnt[0] ),
    .A2(\u_timer.u_pulse_1us.cnt[1] ),
    .B1(\u_timer.u_pulse_1us.cnt[2] ),
    .X(_03935_));
 sky130_fd_sc_hd__and3_1 _08823_ (.A(_01531_),
    .B(_03934_),
    .C(_03935_),
    .X(_00502_));
 sky130_fd_sc_hd__nor2_1 _08824_ (.A(_00928_),
    .B(_03934_),
    .Y(_03936_));
 sky130_fd_sc_hd__o21ai_1 _08825_ (.A1(\u_timer.u_pulse_1us.cnt[3] ),
    .A2(_03933_),
    .B1(_01531_),
    .Y(_03937_));
 sky130_fd_sc_hd__nor2_1 _08826_ (.A(_03936_),
    .B(_03937_),
    .Y(_00503_));
 sky130_fd_sc_hd__and3_1 _08827_ (.A(\u_timer.u_pulse_1us.cnt[3] ),
    .B(\u_timer.u_pulse_1us.cnt[4] ),
    .C(_03933_),
    .X(_03938_));
 sky130_fd_sc_hd__o21ai_1 _08828_ (.A1(\u_timer.u_pulse_1us.cnt[4] ),
    .A2(_03936_),
    .B1(_01531_),
    .Y(_03939_));
 sky130_fd_sc_hd__nor2_1 _08829_ (.A(_03938_),
    .B(_03939_),
    .Y(_00504_));
 sky130_fd_sc_hd__and3_1 _08830_ (.A(\u_timer.u_pulse_1us.cnt[4] ),
    .B(\u_timer.u_pulse_1us.cnt[5] ),
    .C(_03936_),
    .X(_03940_));
 sky130_fd_sc_hd__o21ai_1 _08831_ (.A1(\u_timer.u_pulse_1us.cnt[5] ),
    .A2(_03938_),
    .B1(_01531_),
    .Y(_03941_));
 sky130_fd_sc_hd__nor2_1 _08832_ (.A(_03940_),
    .B(_03941_),
    .Y(_00505_));
 sky130_fd_sc_hd__or2_1 _08833_ (.A(\u_timer.u_pulse_1us.cnt[6] ),
    .B(_03940_),
    .X(_03942_));
 sky130_fd_sc_hd__nand2_1 _08834_ (.A(\u_timer.u_pulse_1us.cnt[6] ),
    .B(_03940_),
    .Y(_03943_));
 sky130_fd_sc_hd__and3_1 _08835_ (.A(_01531_),
    .B(_03942_),
    .C(_03943_),
    .X(_00506_));
 sky130_fd_sc_hd__nand2_1 _08836_ (.A(_00931_),
    .B(_03943_),
    .Y(_03944_));
 sky130_fd_sc_hd__nor2_1 _08837_ (.A(_00931_),
    .B(_03943_),
    .Y(_03945_));
 sky130_fd_sc_hd__inv_2 _08838_ (.A(_03945_),
    .Y(_03946_));
 sky130_fd_sc_hd__and3_1 _08839_ (.A(_01531_),
    .B(_03944_),
    .C(_03946_),
    .X(_00507_));
 sky130_fd_sc_hd__nor2_1 _08840_ (.A(_00933_),
    .B(_03946_),
    .Y(_03947_));
 sky130_fd_sc_hd__o21ai_1 _08841_ (.A1(\u_timer.u_pulse_1us.cnt[8] ),
    .A2(_03945_),
    .B1(_01531_),
    .Y(_03948_));
 sky130_fd_sc_hd__nor2_1 _08842_ (.A(_03947_),
    .B(_03948_),
    .Y(_00508_));
 sky130_fd_sc_hd__or2_1 _08843_ (.A(\u_timer.u_pulse_1us.cnt[9] ),
    .B(_03947_),
    .X(_03949_));
 sky130_fd_sc_hd__o311a_1 _08844_ (.A1(_00933_),
    .A2(_00934_),
    .A3(_03946_),
    .B1(_03949_),
    .C1(_01531_),
    .X(_00509_));
 sky130_fd_sc_hd__mux4_1 _08845_ (.A0(\u_semaphore.reg_0[8] ),
    .A1(\u_semaphore.reg_0[9] ),
    .A2(\u_semaphore.reg_0[10] ),
    .A3(\u_semaphore.reg_0[11] ),
    .S0(net1366),
    .S1(net1357),
    .X(_03950_));
 sky130_fd_sc_hd__or2_1 _08846_ (.A(net1369),
    .B(\u_semaphore.reg_0[14] ),
    .X(_03951_));
 sky130_fd_sc_hd__mux4_2 _08847_ (.A0(\u_semaphore.reg_0[12] ),
    .A1(\u_semaphore.reg_0[13] ),
    .A2(\u_semaphore.reg_0[14] ),
    .A3(\u_semaphore.reg_0[15] ),
    .S0(net1369),
    .S1(net1357),
    .X(_03952_));
 sky130_fd_sc_hd__mux2_1 _08848_ (.A0(_03950_),
    .A1(_03952_),
    .S(net1346),
    .X(_03953_));
 sky130_fd_sc_hd__mux2_1 _08849_ (.A0(\u_semaphore.reg_0[2] ),
    .A1(\u_semaphore.reg_0[3] ),
    .S(net1365),
    .X(_03954_));
 sky130_fd_sc_hd__or2_1 _08850_ (.A(net1275),
    .B(_03954_),
    .X(_03955_));
 sky130_fd_sc_hd__o221a_1 _08851_ (.A1(\u_semaphore.reg_0[1] ),
    .A2(_00999_),
    .B1(net1226),
    .B2(\u_semaphore.reg_0[0] ),
    .C1(_03955_),
    .X(_03956_));
 sky130_fd_sc_hd__mux2_1 _08852_ (.A0(\u_semaphore.reg_0[4] ),
    .A1(\u_semaphore.reg_0[5] ),
    .S(net1365),
    .X(_03957_));
 sky130_fd_sc_hd__mux4_1 _08853_ (.A0(\u_semaphore.reg_0[4] ),
    .A1(\u_semaphore.reg_0[5] ),
    .A2(\u_semaphore.reg_0[6] ),
    .A3(\u_semaphore.reg_0[7] ),
    .S0(net1365),
    .S1(net1359),
    .X(_03958_));
 sky130_fd_sc_hd__o221a_1 _08854_ (.A1(_01130_),
    .A2(_03956_),
    .B1(_03958_),
    .B2(_00997_),
    .C1(_01544_),
    .X(_03959_));
 sky130_fd_sc_hd__o21ai_1 _08855_ (.A1(_00779_),
    .A2(_03953_),
    .B1(_03959_),
    .Y(_03960_));
 sky130_fd_sc_hd__o21a_1 _08856_ (.A1(\u_semaphore.reg_0[0] ),
    .A2(_01544_),
    .B1(_03960_),
    .X(\u_semaphore.reg_out[0] ));
 sky130_fd_sc_hd__mux2_1 _08857_ (.A0(\u_semaphore.reg_0[13] ),
    .A1(\u_semaphore.reg_0[14] ),
    .S(net1369),
    .X(_03961_));
 sky130_fd_sc_hd__a22o_1 _08858_ (.A1(\u_semaphore.reg_0[15] ),
    .A2(net1160),
    .B1(_03961_),
    .B2(net1280),
    .X(_03962_));
 sky130_fd_sc_hd__mux2_1 _08859_ (.A0(\u_semaphore.reg_0[9] ),
    .A1(\u_semaphore.reg_0[10] ),
    .S(net1366),
    .X(_03963_));
 sky130_fd_sc_hd__mux2_1 _08860_ (.A0(\u_semaphore.reg_0[11] ),
    .A1(\u_semaphore.reg_0[12] ),
    .S(net1366),
    .X(_03964_));
 sky130_fd_sc_hd__mux2_1 _08861_ (.A0(_03963_),
    .A1(_03964_),
    .S(net1357),
    .X(_03965_));
 sky130_fd_sc_hd__mux2_1 _08862_ (.A0(_03965_),
    .A1(_03962_),
    .S(net1346),
    .X(_03966_));
 sky130_fd_sc_hd__mux2_1 _08863_ (.A0(\u_semaphore.reg_0[5] ),
    .A1(\u_semaphore.reg_0[6] ),
    .S(net1366),
    .X(_03967_));
 sky130_fd_sc_hd__mux2_1 _08864_ (.A0(\u_semaphore.reg_0[7] ),
    .A1(\u_semaphore.reg_0[8] ),
    .S(net1366),
    .X(_03968_));
 sky130_fd_sc_hd__mux2_1 _08865_ (.A0(_03967_),
    .A1(_03968_),
    .S(net1357),
    .X(_03969_));
 sky130_fd_sc_hd__mux2_1 _08866_ (.A0(\u_semaphore.reg_0[3] ),
    .A1(\u_semaphore.reg_0[4] ),
    .S(net1366),
    .X(_03970_));
 sky130_fd_sc_hd__o21a_1 _08867_ (.A1(\u_semaphore.reg_0[1] ),
    .A2(net1226),
    .B1(net1214),
    .X(_03971_));
 sky130_fd_sc_hd__o221a_1 _08868_ (.A1(\u_semaphore.reg_0[2] ),
    .A2(_00999_),
    .B1(_03970_),
    .B2(net1275),
    .C1(_03971_),
    .X(_03972_));
 sky130_fd_sc_hd__a221o_1 _08869_ (.A1(net1345),
    .A2(_03966_),
    .B1(_03969_),
    .B2(net1182),
    .C1(_03972_),
    .X(_03973_));
 sky130_fd_sc_hd__a21o_1 _08870_ (.A1(\u_semaphore.reg_0[1] ),
    .A2(net1129),
    .B1(_03973_),
    .X(\u_semaphore.reg_out[1] ));
 sky130_fd_sc_hd__o211a_1 _08871_ (.A1(net1264),
    .A2(\u_semaphore.reg_0[15] ),
    .B1(_03951_),
    .C1(net1280),
    .X(_03974_));
 sky130_fd_sc_hd__mux4_1 _08872_ (.A0(\u_semaphore.reg_0[10] ),
    .A1(\u_semaphore.reg_0[11] ),
    .A2(\u_semaphore.reg_0[12] ),
    .A3(\u_semaphore.reg_0[13] ),
    .S0(net1366),
    .S1(net1357),
    .X(_03975_));
 sky130_fd_sc_hd__mux2_1 _08873_ (.A0(_03975_),
    .A1(_03974_),
    .S(net1347),
    .X(_03976_));
 sky130_fd_sc_hd__or2_1 _08874_ (.A(net1358),
    .B(_03954_),
    .X(_03977_));
 sky130_fd_sc_hd__o211a_1 _08875_ (.A1(net1276),
    .A2(_03957_),
    .B1(_03977_),
    .C1(net1214),
    .X(_03978_));
 sky130_fd_sc_hd__mux4_1 _08876_ (.A0(\u_semaphore.reg_0[6] ),
    .A1(\u_semaphore.reg_0[7] ),
    .A2(\u_semaphore.reg_0[8] ),
    .A3(\u_semaphore.reg_0[9] ),
    .S0(net1366),
    .S1(net1357),
    .X(_03979_));
 sky130_fd_sc_hd__a22o_1 _08877_ (.A1(\u_semaphore.reg_0[2] ),
    .A2(net1129),
    .B1(_03979_),
    .B2(net1181),
    .X(_03980_));
 sky130_fd_sc_hd__a211o_1 _08878_ (.A1(net1345),
    .A2(_03976_),
    .B1(_03978_),
    .C1(_03980_),
    .X(\u_semaphore.reg_out[2] ));
 sky130_fd_sc_hd__mux2_1 _08879_ (.A0(_03961_),
    .A1(_03964_),
    .S(net1280),
    .X(_03981_));
 sky130_fd_sc_hd__a21bo_1 _08880_ (.A1(\u_semaphore.reg_0[15] ),
    .A2(net1248),
    .B1_N(net1347),
    .X(_03982_));
 sky130_fd_sc_hd__or2_1 _08881_ (.A(net1347),
    .B(_03981_),
    .X(_03983_));
 sky130_fd_sc_hd__and3_1 _08882_ (.A(net1345),
    .B(_03982_),
    .C(_03983_),
    .X(_03984_));
 sky130_fd_sc_hd__or2_1 _08883_ (.A(net1357),
    .B(_03970_),
    .X(_03985_));
 sky130_fd_sc_hd__o211a_1 _08884_ (.A1(net1275),
    .A2(_03967_),
    .B1(_03985_),
    .C1(net1215),
    .X(_03986_));
 sky130_fd_sc_hd__mux2_1 _08885_ (.A0(_03963_),
    .A1(_03968_),
    .S(net1275),
    .X(_03987_));
 sky130_fd_sc_hd__a22o_1 _08886_ (.A1(\u_semaphore.reg_0[3] ),
    .A2(net1129),
    .B1(_03987_),
    .B2(net1182),
    .X(_03988_));
 sky130_fd_sc_hd__or3_1 _08887_ (.A(_03984_),
    .B(_03986_),
    .C(_03988_),
    .X(\u_semaphore.reg_out[3] ));
 sky130_fd_sc_hd__a22o_1 _08888_ (.A1(\u_semaphore.reg_0[4] ),
    .A2(net1129),
    .B1(_03952_),
    .B2(net1152),
    .X(_03989_));
 sky130_fd_sc_hd__a22o_1 _08889_ (.A1(net1181),
    .A2(_03950_),
    .B1(_03958_),
    .B2(net1215),
    .X(_03990_));
 sky130_fd_sc_hd__or2_1 _08890_ (.A(_03989_),
    .B(_03990_),
    .X(\u_semaphore.reg_out[4] ));
 sky130_fd_sc_hd__a22o_1 _08891_ (.A1(net1153),
    .A2(_03962_),
    .B1(_03969_),
    .B2(net1215),
    .X(_03991_));
 sky130_fd_sc_hd__a22o_1 _08892_ (.A1(\u_semaphore.reg_0[5] ),
    .A2(net1129),
    .B1(_03965_),
    .B2(net1181),
    .X(_03992_));
 sky130_fd_sc_hd__or2_1 _08893_ (.A(_03991_),
    .B(_03992_),
    .X(\u_semaphore.reg_out[5] ));
 sky130_fd_sc_hd__a22o_1 _08894_ (.A1(net1152),
    .A2(_03974_),
    .B1(_03979_),
    .B2(net1215),
    .X(_03993_));
 sky130_fd_sc_hd__a22o_1 _08895_ (.A1(\u_semaphore.reg_0[6] ),
    .A2(net1130),
    .B1(_03975_),
    .B2(net1182),
    .X(_03994_));
 sky130_fd_sc_hd__or2_1 _08896_ (.A(_03993_),
    .B(_03994_),
    .X(\u_semaphore.reg_out[6] ));
 sky130_fd_sc_hd__a22o_1 _08897_ (.A1(\u_semaphore.reg_0[7] ),
    .A2(net1129),
    .B1(_03987_),
    .B2(net1215),
    .X(_03995_));
 sky130_fd_sc_hd__a22o_1 _08898_ (.A1(\u_semaphore.reg_0[15] ),
    .A2(net662),
    .B1(_03981_),
    .B2(net1182),
    .X(_03996_));
 sky130_fd_sc_hd__or2_1 _08899_ (.A(_03995_),
    .B(_03996_),
    .X(\u_semaphore.reg_out[7] ));
 sky130_fd_sc_hd__a22o_1 _08900_ (.A1(\u_semaphore.reg_0[8] ),
    .A2(net1129),
    .B1(_03953_),
    .B2(_00779_),
    .X(\u_semaphore.reg_out[8] ));
 sky130_fd_sc_hd__a22o_1 _08901_ (.A1(\u_semaphore.reg_0[9] ),
    .A2(net1129),
    .B1(_03966_),
    .B2(_00779_),
    .X(\u_semaphore.reg_out[9] ));
 sky130_fd_sc_hd__a22o_1 _08902_ (.A1(\u_semaphore.reg_0[10] ),
    .A2(net1129),
    .B1(_03976_),
    .B2(_00779_),
    .X(\u_semaphore.reg_out[10] ));
 sky130_fd_sc_hd__a32o_1 _08903_ (.A1(_00779_),
    .A2(_03982_),
    .A3(_03983_),
    .B1(\u_semaphore.reg_0[11] ),
    .B2(net1130),
    .X(\u_semaphore.reg_out[11] ));
 sky130_fd_sc_hd__a22o_1 _08904_ (.A1(\u_semaphore.reg_0[12] ),
    .A2(net1130),
    .B1(_03952_),
    .B2(net1215),
    .X(\u_semaphore.reg_out[12] ));
 sky130_fd_sc_hd__a22o_1 _08905_ (.A1(\u_semaphore.reg_0[13] ),
    .A2(net1130),
    .B1(_03962_),
    .B2(net1215),
    .X(\u_semaphore.reg_out[13] ));
 sky130_fd_sc_hd__a22o_1 _08906_ (.A1(\u_semaphore.reg_0[14] ),
    .A2(net1130),
    .B1(_03974_),
    .B2(net1215),
    .X(\u_semaphore.reg_out[14] ));
 sky130_fd_sc_hd__o21a_1 _08907_ (.A1(net1134),
    .A2(net1130),
    .B1(\u_semaphore.reg_0[15] ),
    .X(\u_semaphore.reg_out[15] ));
 sky130_fd_sc_hd__and3_4 _08908_ (.A(net1328),
    .B(\u_pwm.reg_ack_glbl ),
    .C(_01563_),
    .X(_03997_));
 sky130_fd_sc_hd__a21oi_1 _08909_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_oneshot ),
    .A2(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .B1(\u_pwm.u_pwm_0.cfg_pwm_run ),
    .Y(_03998_));
 sky130_fd_sc_hd__a31o_1 _08910_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_run ),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_oneshot ),
    .A3(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .B1(_03997_),
    .X(_03999_));
 sky130_fd_sc_hd__a21oi_1 _08911_ (.A1(net1428),
    .A2(_03997_),
    .B1(\u_pwm.u_pwm_0.gpio_tgr ),
    .Y(_04000_));
 sky130_fd_sc_hd__o21ai_1 _08912_ (.A1(_03998_),
    .A2(_03999_),
    .B1(_04000_),
    .Y(_00308_));
 sky130_fd_sc_hd__a21oi_1 _08913_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_oneshot ),
    .A2(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .B1(\u_pwm.u_pwm_1.cfg_pwm_run ),
    .Y(_04001_));
 sky130_fd_sc_hd__a311oi_1 _08914_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_run ),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_oneshot ),
    .A3(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .B1(_03997_),
    .C1(_04001_),
    .Y(_04002_));
 sky130_fd_sc_hd__a211o_1 _08915_ (.A1(net1421),
    .A2(_03997_),
    .B1(_04002_),
    .C1(\u_pwm.u_pwm_1.gpio_tgr ),
    .X(_00309_));
 sky130_fd_sc_hd__nand2_1 _08916_ (.A(\u_pwm.u_pwm_2.cfg_pwm_oneshot ),
    .B(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .Y(_04003_));
 sky130_fd_sc_hd__xor2_1 _08917_ (.A(\u_pwm.u_pwm_2.cfg_pwm_run ),
    .B(_04003_),
    .X(_04004_));
 sky130_fd_sc_hd__nor2_1 _08918_ (.A(_03997_),
    .B(_04004_),
    .Y(_04005_));
 sky130_fd_sc_hd__a211o_1 _08919_ (.A1(net1289),
    .A2(_03997_),
    .B1(_04005_),
    .C1(\u_pwm.u_pwm_2.gpio_tgr ),
    .X(_00310_));
 sky130_fd_sc_hd__and2_1 _08920_ (.A(_01386_),
    .B(net677),
    .X(_04006_));
 sky130_fd_sc_hd__and3_1 _08921_ (.A(_00873_),
    .B(_01386_),
    .C(net677),
    .X(_00319_));
 sky130_fd_sc_hd__o21ai_1 _08922_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .B1(net513),
    .Y(_04007_));
 sky130_fd_sc_hd__a21oi_1 _08923_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .B1(_04007_),
    .Y(_00326_));
 sky130_fd_sc_hd__a21o_1 _08924_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ),
    .X(_04008_));
 sky130_fd_sc_hd__and3b_1 _08925_ (.A_N(_01356_),
    .B(net514),
    .C(_04008_),
    .X(_00327_));
 sky130_fd_sc_hd__or2_1 _08926_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ),
    .B(_01356_),
    .X(_04009_));
 sky130_fd_sc_hd__and3b_1 _08927_ (.A_N(_01357_),
    .B(net514),
    .C(_04009_),
    .X(_00328_));
 sky130_fd_sc_hd__o21ai_1 _08928_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .A2(_01357_),
    .B1(net514),
    .Y(_04010_));
 sky130_fd_sc_hd__a21oi_1 _08929_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .A2(_01357_),
    .B1(_04010_),
    .Y(_00329_));
 sky130_fd_sc_hd__a21o_1 _08930_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ),
    .A2(_01357_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ),
    .X(_04011_));
 sky130_fd_sc_hd__and3b_1 _08931_ (.A_N(_01358_),
    .B(net514),
    .C(_04011_),
    .X(_00330_));
 sky130_fd_sc_hd__o21ai_1 _08932_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ),
    .A2(_01358_),
    .B1(net514),
    .Y(_04012_));
 sky130_fd_sc_hd__nor2_1 _08933_ (.A(_01359_),
    .B(_04012_),
    .Y(_00331_));
 sky130_fd_sc_hd__o21ai_1 _08934_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ),
    .A2(_01359_),
    .B1(net513),
    .Y(_04013_));
 sky130_fd_sc_hd__nor2_1 _08935_ (.A(_01360_),
    .B(_04013_),
    .Y(_00332_));
 sky130_fd_sc_hd__o21ai_1 _08936_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ),
    .A2(_01360_),
    .B1(net513),
    .Y(_04014_));
 sky130_fd_sc_hd__nor2_1 _08937_ (.A(_01361_),
    .B(_04014_),
    .Y(_00333_));
 sky130_fd_sc_hd__o21ai_1 _08938_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .A2(_01361_),
    .B1(net513),
    .Y(_04015_));
 sky130_fd_sc_hd__nor2_1 _08939_ (.A(_01362_),
    .B(_04015_),
    .Y(_00334_));
 sky130_fd_sc_hd__o21ai_1 _08940_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .A2(_01362_),
    .B1(net513),
    .Y(_04016_));
 sky130_fd_sc_hd__a21oi_1 _08941_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .A2(_01362_),
    .B1(_04016_),
    .Y(_00320_));
 sky130_fd_sc_hd__a31o_1 _08942_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ),
    .A3(_01361_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ),
    .X(_04017_));
 sky130_fd_sc_hd__and3b_1 _08943_ (.A_N(_01363_),
    .B(net513),
    .C(_04017_),
    .X(_00321_));
 sky130_fd_sc_hd__o21ai_1 _08944_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .A2(_01363_),
    .B1(net513),
    .Y(_04018_));
 sky130_fd_sc_hd__nor2_1 _08945_ (.A(_01364_),
    .B(_04018_),
    .Y(_00322_));
 sky130_fd_sc_hd__o21ai_1 _08946_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .A2(_01364_),
    .B1(net513),
    .Y(_04019_));
 sky130_fd_sc_hd__a21oi_1 _08947_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .A2(_01364_),
    .B1(_04019_),
    .Y(_00323_));
 sky130_fd_sc_hd__a31o_1 _08948_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ),
    .A3(_01363_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ),
    .X(_04020_));
 sky130_fd_sc_hd__and3b_1 _08949_ (.A_N(_01365_),
    .B(net513),
    .C(_04020_),
    .X(_00324_));
 sky130_fd_sc_hd__o21a_1 _08950_ (.A1(net1077),
    .A2(_01365_),
    .B1(net513),
    .X(_00325_));
 sky130_fd_sc_hd__and2b_1 _08951_ (.A_N(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ),
    .B(net676),
    .X(_00335_));
 sky130_fd_sc_hd__o21ai_1 _08952_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ),
    .B1(net676),
    .Y(_04021_));
 sky130_fd_sc_hd__nor2_1 _08953_ (.A(_01464_),
    .B(_04021_),
    .Y(_00341_));
 sky130_fd_sc_hd__o21ai_1 _08954_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ),
    .A2(_01464_),
    .B1(net676),
    .Y(_04022_));
 sky130_fd_sc_hd__a21oi_1 _08955_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ),
    .A2(_01464_),
    .B1(_04022_),
    .Y(_00342_));
 sky130_fd_sc_hd__a31o_1 _08956_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ),
    .A2(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ),
    .A3(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[3] ),
    .X(_04023_));
 sky130_fd_sc_hd__and3b_1 _08957_ (.A_N(_01465_),
    .B(_04023_),
    .C(net676),
    .X(_00343_));
 sky130_fd_sc_hd__o21ai_1 _08958_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ),
    .A2(_01465_),
    .B1(net676),
    .Y(_04024_));
 sky130_fd_sc_hd__a21oi_1 _08959_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ),
    .A2(_01465_),
    .B1(_04024_),
    .Y(_00344_));
 sky130_fd_sc_hd__a21o_1 _08960_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ),
    .A2(_01465_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[5] ),
    .X(_04025_));
 sky130_fd_sc_hd__and3b_1 _08961_ (.A_N(_01474_),
    .B(_04025_),
    .C(net676),
    .X(_00345_));
 sky130_fd_sc_hd__o21ai_1 _08962_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ),
    .A2(_01474_),
    .B1(net676),
    .Y(_04026_));
 sky130_fd_sc_hd__a21oi_1 _08963_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ),
    .A2(_01474_),
    .B1(_04026_),
    .Y(_00346_));
 sky130_fd_sc_hd__a21o_1 _08964_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ),
    .A2(_01474_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[7] ),
    .X(_04027_));
 sky130_fd_sc_hd__and3b_1 _08965_ (.A_N(_01475_),
    .B(_04027_),
    .C(net676),
    .X(_00347_));
 sky130_fd_sc_hd__o21ai_1 _08966_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ),
    .A2(_01475_),
    .B1(net676),
    .Y(_04028_));
 sky130_fd_sc_hd__a21oi_1 _08967_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ),
    .A2(_01475_),
    .B1(_04028_),
    .Y(_00348_));
 sky130_fd_sc_hd__a21o_1 _08968_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ),
    .A2(_01475_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[9] ),
    .X(_04029_));
 sky130_fd_sc_hd__and3_1 _08969_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[9] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ),
    .C(_01475_),
    .X(_04030_));
 sky130_fd_sc_hd__and3b_1 _08970_ (.A_N(_04030_),
    .B(net677),
    .C(_04029_),
    .X(_00349_));
 sky130_fd_sc_hd__o21ai_1 _08971_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ),
    .A2(_04030_),
    .B1(net677),
    .Y(_04031_));
 sky130_fd_sc_hd__a21oi_1 _08972_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ),
    .A2(_04030_),
    .B1(_04031_),
    .Y(_00336_));
 sky130_fd_sc_hd__a21o_1 _08973_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ),
    .A2(_04030_),
    .B1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[11] ),
    .X(_04032_));
 sky130_fd_sc_hd__and3_1 _08974_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[11] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ),
    .C(_04030_),
    .X(_04033_));
 sky130_fd_sc_hd__and3b_1 _08975_ (.A_N(_04033_),
    .B(net677),
    .C(_04032_),
    .X(_00337_));
 sky130_fd_sc_hd__and2_1 _08976_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ),
    .B(_04033_),
    .X(_04034_));
 sky130_fd_sc_hd__o21ai_1 _08977_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ),
    .A2(_04033_),
    .B1(net677),
    .Y(_04035_));
 sky130_fd_sc_hd__nor2_1 _08978_ (.A(_04034_),
    .B(_04035_),
    .Y(_00338_));
 sky130_fd_sc_hd__and3_1 _08979_ (.A(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[13] ),
    .B(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ),
    .C(_04033_),
    .X(_04036_));
 sky130_fd_sc_hd__o21ai_1 _08980_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[13] ),
    .A2(_04034_),
    .B1(net677),
    .Y(_04037_));
 sky130_fd_sc_hd__nor2_1 _08981_ (.A(_04036_),
    .B(_04037_),
    .Y(_00339_));
 sky130_fd_sc_hd__a21boi_1 _08982_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[14] ),
    .A2(_04036_),
    .B1_N(net677),
    .Y(_04038_));
 sky130_fd_sc_hd__o21a_1 _08983_ (.A1(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[14] ),
    .A2(_04036_),
    .B1(_04038_),
    .X(_00340_));
 sky130_fd_sc_hd__and2b_1 _08984_ (.A_N(_01426_),
    .B(_01482_),
    .X(_04039_));
 sky130_fd_sc_hd__and2_1 _08985_ (.A(_00893_),
    .B(net518),
    .X(_00372_));
 sky130_fd_sc_hd__or2_1 _08986_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ),
    .X(_04040_));
 sky130_fd_sc_hd__and3_1 _08987_ (.A(_01392_),
    .B(net518),
    .C(_04040_),
    .X(_00379_));
 sky130_fd_sc_hd__nand2_1 _08988_ (.A(_00891_),
    .B(_01392_),
    .Y(_04041_));
 sky130_fd_sc_hd__and3b_1 _08989_ (.A_N(_01393_),
    .B(net518),
    .C(_04041_),
    .X(_00380_));
 sky130_fd_sc_hd__or2_1 _08990_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ),
    .B(_01393_),
    .X(_04042_));
 sky130_fd_sc_hd__and3b_1 _08991_ (.A_N(_01394_),
    .B(net518),
    .C(_04042_),
    .X(_00381_));
 sky130_fd_sc_hd__or2_1 _08992_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ),
    .B(_01394_),
    .X(_04043_));
 sky130_fd_sc_hd__and3_1 _08993_ (.A(_01395_),
    .B(net518),
    .C(_04043_),
    .X(_00382_));
 sky130_fd_sc_hd__nand2_1 _08994_ (.A(net726),
    .B(_01395_),
    .Y(_04044_));
 sky130_fd_sc_hd__and3b_1 _08995_ (.A_N(_01396_),
    .B(net518),
    .C(_04044_),
    .X(_00383_));
 sky130_fd_sc_hd__or2_1 _08996_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ),
    .B(_01396_),
    .X(_04045_));
 sky130_fd_sc_hd__and3b_1 _08997_ (.A_N(_01397_),
    .B(net517),
    .C(_04045_),
    .X(_00384_));
 sky130_fd_sc_hd__or2_1 _08998_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ),
    .B(_01397_),
    .X(_04046_));
 sky130_fd_sc_hd__and3_1 _08999_ (.A(_01398_),
    .B(net517),
    .C(_04046_),
    .X(_00385_));
 sky130_fd_sc_hd__nand2_1 _09000_ (.A(_00885_),
    .B(_01398_),
    .Y(_04047_));
 sky130_fd_sc_hd__and3b_1 _09001_ (.A_N(_01399_),
    .B(net517),
    .C(_04047_),
    .X(_00386_));
 sky130_fd_sc_hd__or2_1 _09002_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ),
    .B(_01399_),
    .X(_04048_));
 sky130_fd_sc_hd__and3b_1 _09003_ (.A_N(_01400_),
    .B(net517),
    .C(_04048_),
    .X(_00387_));
 sky130_fd_sc_hd__or2_1 _09004_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ),
    .B(_01400_),
    .X(_04049_));
 sky130_fd_sc_hd__and3_1 _09005_ (.A(_01401_),
    .B(net517),
    .C(_04049_),
    .X(_00373_));
 sky130_fd_sc_hd__nand2_1 _09006_ (.A(_00882_),
    .B(_01401_),
    .Y(_04050_));
 sky130_fd_sc_hd__and3b_1 _09007_ (.A_N(_01402_),
    .B(net517),
    .C(_04050_),
    .X(_00374_));
 sky130_fd_sc_hd__or2_1 _09008_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ),
    .B(_01402_),
    .X(_04051_));
 sky130_fd_sc_hd__and3b_1 _09009_ (.A_N(_01403_),
    .B(net517),
    .C(_04051_),
    .X(_00375_));
 sky130_fd_sc_hd__or2_1 _09010_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ),
    .B(_01403_),
    .X(_04052_));
 sky130_fd_sc_hd__and3_1 _09011_ (.A(_01404_),
    .B(net517),
    .C(_04052_),
    .X(_00376_));
 sky130_fd_sc_hd__nand2_1 _09012_ (.A(_00879_),
    .B(_01404_),
    .Y(_04053_));
 sky130_fd_sc_hd__and3b_1 _09013_ (.A_N(_01405_),
    .B(net517),
    .C(_04053_),
    .X(_00377_));
 sky130_fd_sc_hd__o21a_1 _09014_ (.A1(net1074),
    .A2(_01405_),
    .B1(net517),
    .X(_00378_));
 sky130_fd_sc_hd__and2b_1 _09015_ (.A_N(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ),
    .B(net675),
    .X(_00388_));
 sky130_fd_sc_hd__o21ai_1 _09016_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ),
    .A2(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ),
    .B1(net674),
    .Y(_04054_));
 sky130_fd_sc_hd__nor2_1 _09017_ (.A(_01483_),
    .B(_04054_),
    .Y(_00394_));
 sky130_fd_sc_hd__o21ai_1 _09018_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ),
    .A2(_01483_),
    .B1(net674),
    .Y(_04055_));
 sky130_fd_sc_hd__a21oi_1 _09019_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ),
    .A2(_01483_),
    .B1(_04055_),
    .Y(_00395_));
 sky130_fd_sc_hd__a31o_1 _09020_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ),
    .A2(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ),
    .A3(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[3] ),
    .X(_04056_));
 sky130_fd_sc_hd__and3b_1 _09021_ (.A_N(_01484_),
    .B(_04056_),
    .C(net675),
    .X(_00396_));
 sky130_fd_sc_hd__o21ai_1 _09022_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ),
    .A2(_01484_),
    .B1(net675),
    .Y(_04057_));
 sky130_fd_sc_hd__a21oi_1 _09023_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ),
    .A2(_01484_),
    .B1(_04057_),
    .Y(_00397_));
 sky130_fd_sc_hd__a21o_1 _09024_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ),
    .A2(_01484_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[5] ),
    .X(_04058_));
 sky130_fd_sc_hd__and3b_1 _09025_ (.A_N(_01499_),
    .B(_04058_),
    .C(net675),
    .X(_00398_));
 sky130_fd_sc_hd__o21ai_1 _09026_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ),
    .A2(_01499_),
    .B1(net675),
    .Y(_04059_));
 sky130_fd_sc_hd__a21oi_1 _09027_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ),
    .A2(_01499_),
    .B1(_04059_),
    .Y(_00399_));
 sky130_fd_sc_hd__a21o_1 _09028_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ),
    .A2(_01499_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[7] ),
    .X(_04060_));
 sky130_fd_sc_hd__and3b_1 _09029_ (.A_N(_01500_),
    .B(_04060_),
    .C(net675),
    .X(_00400_));
 sky130_fd_sc_hd__o21ai_1 _09030_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ),
    .A2(_01500_),
    .B1(net674),
    .Y(_04061_));
 sky130_fd_sc_hd__a21oi_1 _09031_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ),
    .A2(_01500_),
    .B1(_04061_),
    .Y(_00401_));
 sky130_fd_sc_hd__a21o_1 _09032_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ),
    .A2(_01500_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[9] ),
    .X(_04062_));
 sky130_fd_sc_hd__and3_1 _09033_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[9] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ),
    .C(_01500_),
    .X(_04063_));
 sky130_fd_sc_hd__and3b_1 _09034_ (.A_N(_04063_),
    .B(net674),
    .C(_04062_),
    .X(_00402_));
 sky130_fd_sc_hd__o21ai_1 _09035_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ),
    .A2(_04063_),
    .B1(net674),
    .Y(_04064_));
 sky130_fd_sc_hd__a21oi_1 _09036_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ),
    .A2(_04063_),
    .B1(_04064_),
    .Y(_00389_));
 sky130_fd_sc_hd__a21o_1 _09037_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ),
    .A2(_04063_),
    .B1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[11] ),
    .X(_04065_));
 sky130_fd_sc_hd__and3_1 _09038_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[11] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ),
    .C(_04063_),
    .X(_04066_));
 sky130_fd_sc_hd__and3b_1 _09039_ (.A_N(_04066_),
    .B(net674),
    .C(_04065_),
    .X(_00390_));
 sky130_fd_sc_hd__and2_1 _09040_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ),
    .B(_04066_),
    .X(_04067_));
 sky130_fd_sc_hd__o21ai_1 _09041_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ),
    .A2(_04066_),
    .B1(net674),
    .Y(_04068_));
 sky130_fd_sc_hd__nor2_1 _09042_ (.A(_04067_),
    .B(_04068_),
    .Y(_00391_));
 sky130_fd_sc_hd__and3_1 _09043_ (.A(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[13] ),
    .B(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ),
    .C(_04066_),
    .X(_04069_));
 sky130_fd_sc_hd__o21ai_1 _09044_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[13] ),
    .A2(_04067_),
    .B1(net674),
    .Y(_04070_));
 sky130_fd_sc_hd__nor2_1 _09045_ (.A(_04069_),
    .B(_04070_),
    .Y(_00392_));
 sky130_fd_sc_hd__a21boi_1 _09046_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[14] ),
    .A2(_04069_),
    .B1_N(net674),
    .Y(_04071_));
 sky130_fd_sc_hd__o21a_1 _09047_ (.A1(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[14] ),
    .A2(_04069_),
    .B1(_04071_),
    .X(_00393_));
 sky130_fd_sc_hd__and2b_1 _09048_ (.A_N(_01460_),
    .B(net672),
    .X(_04072_));
 sky130_fd_sc_hd__and2_1 _09049_ (.A(_00913_),
    .B(net524),
    .X(_00425_));
 sky130_fd_sc_hd__or2_1 _09050_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ),
    .X(_04073_));
 sky130_fd_sc_hd__and3_1 _09051_ (.A(_01429_),
    .B(net524),
    .C(_04073_),
    .X(_00432_));
 sky130_fd_sc_hd__nand2_1 _09052_ (.A(net725),
    .B(_01429_),
    .Y(_04074_));
 sky130_fd_sc_hd__and3b_1 _09053_ (.A_N(_01430_),
    .B(net524),
    .C(_04074_),
    .X(_00433_));
 sky130_fd_sc_hd__or2_1 _09054_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ),
    .B(_01430_),
    .X(_04075_));
 sky130_fd_sc_hd__and3b_1 _09055_ (.A_N(_01431_),
    .B(net524),
    .C(_04075_),
    .X(_00434_));
 sky130_fd_sc_hd__o21ai_1 _09056_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .A2(_01431_),
    .B1(net524),
    .Y(_04076_));
 sky130_fd_sc_hd__a21oi_1 _09057_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .A2(_01431_),
    .B1(_04076_),
    .Y(_00435_));
 sky130_fd_sc_hd__a21o_1 _09058_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ),
    .A2(_01431_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ),
    .X(_04077_));
 sky130_fd_sc_hd__and3b_1 _09059_ (.A_N(_01432_),
    .B(net524),
    .C(_04077_),
    .X(_00436_));
 sky130_fd_sc_hd__o21ai_1 _09060_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ),
    .A2(_01432_),
    .B1(net523),
    .Y(_04078_));
 sky130_fd_sc_hd__nor2_1 _09061_ (.A(_01433_),
    .B(_04078_),
    .Y(_00437_));
 sky130_fd_sc_hd__o21ai_1 _09062_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ),
    .A2(_01433_),
    .B1(net523),
    .Y(_04079_));
 sky130_fd_sc_hd__nor2_1 _09063_ (.A(_01434_),
    .B(_04079_),
    .Y(_00438_));
 sky130_fd_sc_hd__o21ai_1 _09064_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ),
    .A2(_01434_),
    .B1(net523),
    .Y(_04080_));
 sky130_fd_sc_hd__nor2_1 _09065_ (.A(_01435_),
    .B(_04080_),
    .Y(_00439_));
 sky130_fd_sc_hd__o21ai_1 _09066_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .A2(_01435_),
    .B1(net523),
    .Y(_04081_));
 sky130_fd_sc_hd__nor2_1 _09067_ (.A(_01436_),
    .B(_04081_),
    .Y(_00440_));
 sky130_fd_sc_hd__o21ai_1 _09068_ (.A1(net1073),
    .A2(_01436_),
    .B1(net523),
    .Y(_04082_));
 sky130_fd_sc_hd__a21oi_1 _09069_ (.A1(net1073),
    .A2(_01436_),
    .B1(_04082_),
    .Y(_00426_));
 sky130_fd_sc_hd__a31o_1 _09070_ (.A1(net1073),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ),
    .A3(_01435_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ),
    .X(_04083_));
 sky130_fd_sc_hd__and3b_1 _09071_ (.A_N(_01437_),
    .B(net523),
    .C(_04083_),
    .X(_00427_));
 sky130_fd_sc_hd__o21ai_1 _09072_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ),
    .A2(_01437_),
    .B1(net523),
    .Y(_04084_));
 sky130_fd_sc_hd__nor2_1 _09073_ (.A(_01438_),
    .B(_04084_),
    .Y(_00428_));
 sky130_fd_sc_hd__o21ai_1 _09074_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ),
    .A2(_01438_),
    .B1(net523),
    .Y(_04085_));
 sky130_fd_sc_hd__nor2_1 _09075_ (.A(_01439_),
    .B(_04085_),
    .Y(_00429_));
 sky130_fd_sc_hd__o21ai_1 _09076_ (.A1(net1072),
    .A2(_01439_),
    .B1(net523),
    .Y(_04086_));
 sky130_fd_sc_hd__a21oi_1 _09077_ (.A1(net1072),
    .A2(_01439_),
    .B1(_04086_),
    .Y(_00430_));
 sky130_fd_sc_hd__a21o_1 _09078_ (.A1(net1072),
    .A2(_01439_),
    .B1(net1070),
    .X(_04087_));
 sky130_fd_sc_hd__and2_1 _09079_ (.A(net523),
    .B(_04087_),
    .X(_00431_));
 sky130_fd_sc_hd__and2b_1 _09080_ (.A_N(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ),
    .B(net673),
    .X(_00441_));
 sky130_fd_sc_hd__o21ai_1 _09081_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ),
    .B1(net673),
    .Y(_04088_));
 sky130_fd_sc_hd__nor2_1 _09082_ (.A(_01502_),
    .B(_04088_),
    .Y(_00447_));
 sky130_fd_sc_hd__o21ai_1 _09083_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ),
    .A2(_01502_),
    .B1(net673),
    .Y(_04089_));
 sky130_fd_sc_hd__a21oi_1 _09084_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ),
    .A2(_01502_),
    .B1(_04089_),
    .Y(_00448_));
 sky130_fd_sc_hd__a31o_1 _09085_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ),
    .A2(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ),
    .A3(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[3] ),
    .X(_04090_));
 sky130_fd_sc_hd__and3b_1 _09086_ (.A_N(_01503_),
    .B(_04090_),
    .C(net673),
    .X(_00449_));
 sky130_fd_sc_hd__o21ai_1 _09087_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ),
    .A2(_01503_),
    .B1(net673),
    .Y(_04091_));
 sky130_fd_sc_hd__a21oi_1 _09088_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ),
    .A2(_01503_),
    .B1(_04091_),
    .Y(_00450_));
 sky130_fd_sc_hd__a21o_1 _09089_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ),
    .A2(_01503_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[5] ),
    .X(_04092_));
 sky130_fd_sc_hd__and3b_1 _09090_ (.A_N(_01512_),
    .B(_04092_),
    .C(net673),
    .X(_00451_));
 sky130_fd_sc_hd__o21ai_1 _09091_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ),
    .A2(_01512_),
    .B1(net672),
    .Y(_04093_));
 sky130_fd_sc_hd__a21oi_1 _09092_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ),
    .A2(_01512_),
    .B1(_04093_),
    .Y(_00452_));
 sky130_fd_sc_hd__a21o_1 _09093_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ),
    .A2(_01512_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[7] ),
    .X(_04094_));
 sky130_fd_sc_hd__and3b_1 _09094_ (.A_N(_01513_),
    .B(_04094_),
    .C(net672),
    .X(_00453_));
 sky130_fd_sc_hd__o21ai_1 _09095_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ),
    .A2(_01513_),
    .B1(net672),
    .Y(_04095_));
 sky130_fd_sc_hd__a21oi_1 _09096_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ),
    .A2(_01513_),
    .B1(_04095_),
    .Y(_00454_));
 sky130_fd_sc_hd__a21o_1 _09097_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ),
    .A2(_01513_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[9] ),
    .X(_04096_));
 sky130_fd_sc_hd__and3_1 _09098_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[9] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ),
    .C(_01513_),
    .X(_04097_));
 sky130_fd_sc_hd__and3b_1 _09099_ (.A_N(_04097_),
    .B(net672),
    .C(_04096_),
    .X(_00455_));
 sky130_fd_sc_hd__o21ai_1 _09100_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ),
    .A2(_04097_),
    .B1(net672),
    .Y(_04098_));
 sky130_fd_sc_hd__a21oi_1 _09101_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ),
    .A2(_04097_),
    .B1(_04098_),
    .Y(_00442_));
 sky130_fd_sc_hd__a21o_1 _09102_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ),
    .A2(_04097_),
    .B1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[11] ),
    .X(_04099_));
 sky130_fd_sc_hd__and3_1 _09103_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[11] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ),
    .C(_04097_),
    .X(_04100_));
 sky130_fd_sc_hd__and3b_1 _09104_ (.A_N(_04100_),
    .B(net673),
    .C(_04099_),
    .X(_00443_));
 sky130_fd_sc_hd__and2_1 _09105_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ),
    .B(_04100_),
    .X(_04101_));
 sky130_fd_sc_hd__o21ai_1 _09106_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ),
    .A2(_04100_),
    .B1(net672),
    .Y(_04102_));
 sky130_fd_sc_hd__nor2_1 _09107_ (.A(_04101_),
    .B(_04102_),
    .Y(_00444_));
 sky130_fd_sc_hd__and3_1 _09108_ (.A(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[13] ),
    .B(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ),
    .C(_04100_),
    .X(_04103_));
 sky130_fd_sc_hd__o21ai_1 _09109_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[13] ),
    .A2(_04101_),
    .B1(net672),
    .Y(_04104_));
 sky130_fd_sc_hd__nor2_1 _09110_ (.A(_04103_),
    .B(_04104_),
    .Y(_00445_));
 sky130_fd_sc_hd__a21boi_1 _09111_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[14] ),
    .A2(_04103_),
    .B1_N(net672),
    .Y(_04105_));
 sky130_fd_sc_hd__o21a_1 _09112_ (.A1(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[14] ),
    .A2(_04103_),
    .B1(_04105_),
    .X(_00446_));
 sky130_fd_sc_hd__and2_4 _09113_ (.A(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .B(net22),
    .X(net329));
 sky130_fd_sc_hd__and2_4 _09114_ (.A(\u_glbl_reg.cfg_multi_func_sel[15] ),
    .B(net21),
    .X(net330));
 sky130_fd_sc_hd__and2_2 _09115_ (.A(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .B(net1417),
    .X(net460));
 sky130_fd_sc_hd__and2_2 _09116_ (.A(\u_glbl_reg.cfg_multi_func_sel[9] ),
    .B(net1387),
    .X(net502));
 sky130_fd_sc_hd__or3b_1 _09117_ (.A(net1388),
    .B(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .C_N(\u_glbl_reg.cfg_multi_func_sel[8] ),
    .X(net501));
 sky130_fd_sc_hd__and2_4 _09118_ (.A(\u_gpio.cfg_gpio_out_data[17] ),
    .B(\u_gpio.cfg_gpio_dir_sel[17] ),
    .X(net306));
 sky130_fd_sc_hd__and2_4 _09119_ (.A(\u_gpio.cfg_gpio_out_data[16] ),
    .B(\u_gpio.cfg_gpio_dir_sel[16] ),
    .X(net305));
 sky130_fd_sc_hd__o21bai_4 _09120_ (.A1(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[3] ),
    .B1_N(net1109),
    .Y(net284));
 sky130_fd_sc_hd__o21bai_4 _09121_ (.A1(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[2] ),
    .B1_N(net1109),
    .Y(net275));
 sky130_fd_sc_hd__o21bai_4 _09122_ (.A1(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[1] ),
    .B1_N(net1109),
    .Y(net264));
 sky130_fd_sc_hd__o21bai_4 _09123_ (.A1(\u_glbl_reg.cfg_multi_func_sel[18] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[0] ),
    .B1_N(\u_glbl_reg.cfg_multi_func_sel[30] ),
    .Y(net253));
 sky130_fd_sc_hd__or2_1 _09124_ (.A(net1652),
    .B(net1406),
    .X(net282));
 sky130_fd_sc_hd__or2_1 _09125_ (.A(net1652),
    .B(net1408),
    .X(net281));
 sky130_fd_sc_hd__or2_1 _09126_ (.A(net1652),
    .B(net1410),
    .X(net280));
 sky130_fd_sc_hd__or2_1 _09127_ (.A(net1652),
    .B(net1412),
    .X(net279));
 sky130_fd_sc_hd__o31ai_4 _09128_ (.A1(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .A2(\u_gpio.cfg_gpio_dir_sel[12] ),
    .A3(\u_gpio.cfg_gpio_out_type[12] ),
    .B1(_00987_),
    .Y(net265));
 sky130_fd_sc_hd__or4b_1 _09129_ (.A(\u_glbl_reg.cfg_multi_func_sel[5] ),
    .B(\u_gpio.cfg_gpio_dir_sel[11] ),
    .C(\u_gpio.cfg_gpio_out_type[11] ),
    .D_N(net34),
    .X(_04106_));
 sky130_fd_sc_hd__or3b_4 _09130_ (.A(\u_glbl_reg.cfg_multi_func_sel[10] ),
    .B(net1651),
    .C_N(_04106_),
    .X(net263));
 sky130_fd_sc_hd__or4_2 _09131_ (.A(\u_glbl_reg.cfg_multi_func_sel[4] ),
    .B(\u_gpio.cfg_gpio_dir_sel[10] ),
    .C(\u_gpio.cfg_gpio_out_type[10] ),
    .D(\u_glbl_reg.cfg_multi_func_sel[11] ),
    .X(_04107_));
 sky130_fd_sc_hd__nand2_1 _09132_ (.A(_00987_),
    .B(_04107_),
    .Y(net262));
 sky130_fd_sc_hd__or4_2 _09133_ (.A(\u_glbl_reg.cfg_multi_func_sel[3] ),
    .B(\u_gpio.cfg_gpio_dir_sel[9] ),
    .C(\u_gpio.cfg_gpio_out_type[9] ),
    .D(\u_glbl_reg.cfg_multi_func_sel[12] ),
    .X(_04108_));
 sky130_fd_sc_hd__nand2_1 _09134_ (.A(_00987_),
    .B(_04108_),
    .Y(net261));
 sky130_fd_sc_hd__o21ai_2 _09135_ (.A1(\u_gpio.cfg_gpio_dir_sel[8] ),
    .A2(\u_gpio.cfg_gpio_out_type[8] ),
    .B1(_00987_),
    .Y(net260));
 sky130_fd_sc_hd__o31ai_2 _09136_ (.A1(\u_gpio.cfg_gpio_dir_sel[31] ),
    .A2(\u_gpio.cfg_gpio_out_type[31] ),
    .A3(\u_glbl_reg.cfg_multi_func_sel[17] ),
    .B1(_00987_),
    .Y(net259));
 sky130_fd_sc_hd__or4_4 _09137_ (.A(\u_gpio.cfg_gpio_dir_sel[30] ),
    .B(\u_gpio.cfg_gpio_out_type[30] ),
    .C(\u_glbl_reg.cfg_multi_func_sel[13] ),
    .D(\u_glbl_reg.cfg_multi_func_sel[2] ),
    .X(_04109_));
 sky130_fd_sc_hd__nand2_2 _09138_ (.A(_00987_),
    .B(_04109_),
    .Y(net258));
 sky130_fd_sc_hd__or4_2 _09139_ (.A(\u_gpio.cfg_gpio_dir_sel[29] ),
    .B(\u_gpio.cfg_gpio_out_type[29] ),
    .C(\u_glbl_reg.cfg_multi_func_sel[14] ),
    .D(\u_glbl_reg.cfg_multi_func_sel[1] ),
    .X(_04110_));
 sky130_fd_sc_hd__nand2_2 _09140_ (.A(_00987_),
    .B(_04110_),
    .Y(net257));
 sky130_fd_sc_hd__o21bai_4 _09141_ (.A1(\u_gpio.cfg_gpio_dir_sel[26] ),
    .A2(\u_gpio.cfg_gpio_out_type[26] ),
    .B1_N(\u_glbl_reg.cfg_multi_func_sel[6] ),
    .Y(net289));
 sky130_fd_sc_hd__or3_4 _09142_ (.A(\u_glbl_reg.cfg_multi_func_sel[31] ),
    .B(\u_glbl_reg.cfg_multi_func_sel[8] ),
    .C(_01611_),
    .X(net287));
 sky130_fd_sc_hd__nor2_1 _09143_ (.A(_00988_),
    .B(net463),
    .Y(net461));
 sky130_fd_sc_hd__and2_4 _09144_ (.A(net1109),
    .B(net14),
    .X(net450));
 sky130_fd_sc_hd__and2_2 _09145_ (.A(net1109),
    .B(net24),
    .X(net452));
 sky130_fd_sc_hd__and2_4 _09146_ (.A(net1109),
    .B(net32),
    .X(net451));
 sky130_fd_sc_hd__o21ai_1 _09147_ (.A1(\u_glbl_reg.dbg_clk_div16 ),
    .A2(_01108_),
    .B1(_00045_),
    .Y(_00043_));
 sky130_fd_sc_hd__o21ai_1 _09148_ (.A1(net365),
    .A2(_01112_),
    .B1(_00055_),
    .Y(_00053_));
 sky130_fd_sc_hd__xor2_4 _09149_ (.A(\u_glbl_reg.u_random.s1[0] ),
    .B(\u_glbl_reg.u_random.s0[0] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[0] ));
 sky130_fd_sc_hd__xor2_1 _09150_ (.A(\u_glbl_reg.u_random.s0[6] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[0] ),
    .X(_00023_));
 sky130_fd_sc_hd__xor2_4 _09151_ (.A(\u_glbl_reg.u_random.s1[1] ),
    .B(\u_glbl_reg.u_random.s0[1] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[1] ));
 sky130_fd_sc_hd__xor2_1 _09152_ (.A(\u_glbl_reg.u_random.s0[7] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[1] ),
    .X(_00024_));
 sky130_fd_sc_hd__xor2_2 _09153_ (.A(\u_glbl_reg.u_random.s1[2] ),
    .B(\u_glbl_reg.u_random.s0[2] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[2] ));
 sky130_fd_sc_hd__xor2_1 _09154_ (.A(\u_glbl_reg.u_random.s0[8] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[2] ),
    .X(_00025_));
 sky130_fd_sc_hd__xor2_2 _09155_ (.A(\u_glbl_reg.u_random.s1[3] ),
    .B(\u_glbl_reg.u_random.s0[3] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[3] ));
 sky130_fd_sc_hd__xor2_1 _09156_ (.A(\u_glbl_reg.u_random.s0[9] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[3] ),
    .X(_00026_));
 sky130_fd_sc_hd__xor2_2 _09157_ (.A(\u_glbl_reg.u_random.s1[4] ),
    .B(\u_glbl_reg.u_random.s0[4] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[4] ));
 sky130_fd_sc_hd__xor2_1 _09158_ (.A(\u_glbl_reg.u_random.s0[10] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[4] ),
    .X(_00027_));
 sky130_fd_sc_hd__xor2_2 _09159_ (.A(\u_glbl_reg.u_random.s1[5] ),
    .B(\u_glbl_reg.u_random.s0[5] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[5] ));
 sky130_fd_sc_hd__xor2_1 _09160_ (.A(\u_glbl_reg.u_random.s0[11] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[5] ),
    .X(_00028_));
 sky130_fd_sc_hd__xor2_4 _09161_ (.A(\u_glbl_reg.u_random.s0[6] ),
    .B(\u_glbl_reg.u_random.s1[6] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[6] ));
 sky130_fd_sc_hd__xor2_1 _09162_ (.A(\u_glbl_reg.u_random.s0[12] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[6] ),
    .X(_00029_));
 sky130_fd_sc_hd__xor2_2 _09163_ (.A(\u_glbl_reg.u_random.s0[7] ),
    .B(\u_glbl_reg.u_random.s1[7] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[7] ));
 sky130_fd_sc_hd__xor2_1 _09164_ (.A(\u_glbl_reg.u_random.s0[13] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[7] ),
    .X(_00030_));
 sky130_fd_sc_hd__xor2_2 _09165_ (.A(\u_glbl_reg.u_random.s0[8] ),
    .B(\u_glbl_reg.u_random.s1[8] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[8] ));
 sky130_fd_sc_hd__xor2_1 _09166_ (.A(\u_glbl_reg.u_random.s0[14] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[8] ),
    .X(_00031_));
 sky130_fd_sc_hd__xor2_2 _09167_ (.A(\u_glbl_reg.u_random.s0[9] ),
    .B(\u_glbl_reg.u_random.s1[9] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[9] ));
 sky130_fd_sc_hd__xor2_2 _09168_ (.A(\u_glbl_reg.u_random.s0[10] ),
    .B(\u_glbl_reg.u_random.s1[10] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[10] ));
 sky130_fd_sc_hd__xor2_2 _09169_ (.A(\u_glbl_reg.u_random.s0[11] ),
    .B(\u_glbl_reg.u_random.s1[11] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[11] ));
 sky130_fd_sc_hd__xor2_2 _09170_ (.A(\u_glbl_reg.u_random.s0[12] ),
    .B(\u_glbl_reg.u_random.s1[12] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[12] ));
 sky130_fd_sc_hd__xor2_2 _09171_ (.A(\u_glbl_reg.u_random.s0[13] ),
    .B(\u_glbl_reg.u_random.s1[13] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[13] ));
 sky130_fd_sc_hd__xor2_2 _09172_ (.A(\u_glbl_reg.u_random.s0[14] ),
    .B(\u_glbl_reg.u_random.s1[14] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[14] ));
 sky130_fd_sc_hd__xor2_2 _09173_ (.A(\u_glbl_reg.u_random.s1[15] ),
    .B(\u_glbl_reg.u_random.s0[15] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[15] ));
 sky130_fd_sc_hd__xor2_2 _09174_ (.A(\u_glbl_reg.u_random.s1[16] ),
    .B(\u_glbl_reg.u_random.s0[16] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[16] ));
 sky130_fd_sc_hd__xor2_4 _09175_ (.A(\u_glbl_reg.u_random.s1[17] ),
    .B(\u_glbl_reg.u_random.s0[17] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[17] ));
 sky130_fd_sc_hd__xor2_4 _09176_ (.A(\u_glbl_reg.u_random.s1[18] ),
    .B(\u_glbl_reg.u_random.s0[18] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[18] ));
 sky130_fd_sc_hd__xor2_4 _09177_ (.A(\u_glbl_reg.u_random.s1[19] ),
    .B(\u_glbl_reg.u_random.s0[19] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[19] ));
 sky130_fd_sc_hd__xor2_2 _09178_ (.A(\u_glbl_reg.u_random.s1[20] ),
    .B(\u_glbl_reg.u_random.s0[20] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[20] ));
 sky130_fd_sc_hd__xor2_2 _09179_ (.A(\u_glbl_reg.u_random.s1[21] ),
    .B(\u_glbl_reg.u_random.s0[21] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[21] ));
 sky130_fd_sc_hd__xor2_2 _09180_ (.A(\u_glbl_reg.u_random.s1[22] ),
    .B(\u_glbl_reg.u_random.s0[22] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[22] ));
 sky130_fd_sc_hd__xor2_1 _09181_ (.A(\u_glbl_reg.u_random.s1[23] ),
    .B(\u_glbl_reg.u_random.s0[23] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[23] ));
 sky130_fd_sc_hd__xor2_1 _09182_ (.A(\u_glbl_reg.u_random.s1[24] ),
    .B(\u_glbl_reg.u_random.s0[24] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[24] ));
 sky130_fd_sc_hd__xor2_1 _09183_ (.A(\u_glbl_reg.u_random.s1[25] ),
    .B(\u_glbl_reg.u_random.s0[25] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[25] ));
 sky130_fd_sc_hd__xor2_1 _09184_ (.A(\u_glbl_reg.u_random.s1[26] ),
    .B(\u_glbl_reg.u_random.s0[26] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[26] ));
 sky130_fd_sc_hd__xor2_1 _09185_ (.A(\u_glbl_reg.u_random.s1[27] ),
    .B(\u_glbl_reg.u_random.s0[27] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[27] ));
 sky130_fd_sc_hd__xor2_1 _09186_ (.A(\u_glbl_reg.u_random.s1[28] ),
    .B(\u_glbl_reg.u_random.s0[28] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[28] ));
 sky130_fd_sc_hd__xor2_1 _09187_ (.A(\u_glbl_reg.u_random.s1[29] ),
    .B(\u_glbl_reg.u_random.s0[29] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[29] ));
 sky130_fd_sc_hd__xor2_1 _09188_ (.A(\u_glbl_reg.u_random.s1[30] ),
    .B(\u_glbl_reg.u_random.s0[30] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[30] ));
 sky130_fd_sc_hd__xor2_1 _09189_ (.A(\u_glbl_reg.u_random.s1[31] ),
    .B(\u_glbl_reg.u_random.s0[31] ),
    .X(\u_glbl_reg.u_random.s1_xor_s0[31] ));
 sky130_fd_sc_hd__o21ai_1 _09190_ (.A1(\u_glbl_reg.rtc_clk_div ),
    .A2(_01143_),
    .B1(_00194_),
    .Y(_00192_));
 sky130_fd_sc_hd__and2_1 _09191_ (.A(net1474),
    .B(net735),
    .X(_00775_));
 sky130_fd_sc_hd__and3_1 _09192_ (.A(net1474),
    .B(net737),
    .C(net1044),
    .X(_00224_));
 sky130_fd_sc_hd__xnor2_1 _09193_ (.A(\u_glbl_reg.u_random.s0[15] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[9] ),
    .Y(_04111_));
 sky130_fd_sc_hd__xnor2_1 _09194_ (.A(\u_glbl_reg.u_random.s1_xor_s0[0] ),
    .B(_04111_),
    .Y(_00000_));
 sky130_fd_sc_hd__xnor2_1 _09195_ (.A(\u_glbl_reg.u_random.s0[16] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[10] ),
    .Y(_04112_));
 sky130_fd_sc_hd__xnor2_1 _09196_ (.A(\u_glbl_reg.u_random.s1_xor_s0[1] ),
    .B(_04112_),
    .Y(_00011_));
 sky130_fd_sc_hd__xnor2_1 _09197_ (.A(\u_glbl_reg.u_random.s0[17] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[11] ),
    .Y(_04113_));
 sky130_fd_sc_hd__xnor2_1 _09198_ (.A(\u_glbl_reg.u_random.s1_xor_s0[2] ),
    .B(_04113_),
    .Y(_00015_));
 sky130_fd_sc_hd__xnor2_1 _09199_ (.A(\u_glbl_reg.u_random.s0[18] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[12] ),
    .Y(_04114_));
 sky130_fd_sc_hd__xnor2_1 _09200_ (.A(\u_glbl_reg.u_random.s1_xor_s0[3] ),
    .B(_04114_),
    .Y(_00016_));
 sky130_fd_sc_hd__xnor2_1 _09201_ (.A(\u_glbl_reg.u_random.s0[19] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[13] ),
    .Y(_04115_));
 sky130_fd_sc_hd__xnor2_1 _09202_ (.A(\u_glbl_reg.u_random.s1_xor_s0[4] ),
    .B(_04115_),
    .Y(_00017_));
 sky130_fd_sc_hd__xnor2_1 _09203_ (.A(\u_glbl_reg.u_random.s0[20] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[14] ),
    .Y(_04116_));
 sky130_fd_sc_hd__xnor2_1 _09204_ (.A(\u_glbl_reg.u_random.s1_xor_s0[5] ),
    .B(_04116_),
    .Y(_00018_));
 sky130_fd_sc_hd__xnor2_1 _09205_ (.A(\u_glbl_reg.u_random.s0[21] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[15] ),
    .Y(_04117_));
 sky130_fd_sc_hd__xnor2_1 _09206_ (.A(\u_glbl_reg.u_random.s1_xor_s0[6] ),
    .B(_04117_),
    .Y(_00019_));
 sky130_fd_sc_hd__xnor2_1 _09207_ (.A(\u_glbl_reg.u_random.s0[22] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[16] ),
    .Y(_04118_));
 sky130_fd_sc_hd__xnor2_1 _09208_ (.A(\u_glbl_reg.u_random.s1_xor_s0[7] ),
    .B(_04118_),
    .Y(_00020_));
 sky130_fd_sc_hd__xnor2_1 _09209_ (.A(\u_glbl_reg.u_random.s0[23] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[17] ),
    .Y(_04119_));
 sky130_fd_sc_hd__xnor2_1 _09210_ (.A(\u_glbl_reg.u_random.s1_xor_s0[8] ),
    .B(_04119_),
    .Y(_00021_));
 sky130_fd_sc_hd__xnor2_1 _09211_ (.A(\u_glbl_reg.u_random.s0[24] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[18] ),
    .Y(_04120_));
 sky130_fd_sc_hd__xnor2_1 _09212_ (.A(\u_glbl_reg.u_random.s1_xor_s0[9] ),
    .B(_04120_),
    .Y(_00022_));
 sky130_fd_sc_hd__xnor2_1 _09213_ (.A(\u_glbl_reg.u_random.s0[25] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[19] ),
    .Y(_04121_));
 sky130_fd_sc_hd__xnor2_1 _09214_ (.A(\u_glbl_reg.u_random.s1_xor_s0[10] ),
    .B(_04121_),
    .Y(_00001_));
 sky130_fd_sc_hd__xnor2_1 _09215_ (.A(\u_glbl_reg.u_random.s0[26] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[20] ),
    .Y(_04122_));
 sky130_fd_sc_hd__xnor2_1 _09216_ (.A(\u_glbl_reg.u_random.s1_xor_s0[11] ),
    .B(_04122_),
    .Y(_00002_));
 sky130_fd_sc_hd__xnor2_1 _09217_ (.A(\u_glbl_reg.u_random.s0[27] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[21] ),
    .Y(_04123_));
 sky130_fd_sc_hd__xnor2_1 _09218_ (.A(\u_glbl_reg.u_random.s1_xor_s0[12] ),
    .B(_04123_),
    .Y(_00003_));
 sky130_fd_sc_hd__xnor2_1 _09219_ (.A(\u_glbl_reg.u_random.s0[28] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[22] ),
    .Y(_04124_));
 sky130_fd_sc_hd__xnor2_1 _09220_ (.A(\u_glbl_reg.u_random.s1_xor_s0[13] ),
    .B(_04124_),
    .Y(_00004_));
 sky130_fd_sc_hd__xnor2_1 _09221_ (.A(\u_glbl_reg.u_random.s0[29] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[23] ),
    .Y(_04125_));
 sky130_fd_sc_hd__xnor2_1 _09222_ (.A(\u_glbl_reg.u_random.s1_xor_s0[14] ),
    .B(_04125_),
    .Y(_00005_));
 sky130_fd_sc_hd__xnor2_1 _09223_ (.A(\u_glbl_reg.u_random.s0[30] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[24] ),
    .Y(_04126_));
 sky130_fd_sc_hd__xnor2_1 _09224_ (.A(\u_glbl_reg.u_random.s1_xor_s0[15] ),
    .B(_04126_),
    .Y(_00006_));
 sky130_fd_sc_hd__xnor2_1 _09225_ (.A(\u_glbl_reg.u_random.s0[31] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[25] ),
    .Y(_04127_));
 sky130_fd_sc_hd__xnor2_1 _09226_ (.A(\u_glbl_reg.u_random.s1_xor_s0[16] ),
    .B(_04127_),
    .Y(_00007_));
 sky130_fd_sc_hd__xnor2_1 _09227_ (.A(\u_glbl_reg.u_random.s0[0] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[26] ),
    .Y(_04128_));
 sky130_fd_sc_hd__xnor2_1 _09228_ (.A(\u_glbl_reg.u_random.s1_xor_s0[17] ),
    .B(_04128_),
    .Y(_00008_));
 sky130_fd_sc_hd__xnor2_1 _09229_ (.A(\u_glbl_reg.u_random.s0[1] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[27] ),
    .Y(_04129_));
 sky130_fd_sc_hd__xnor2_1 _09230_ (.A(\u_glbl_reg.u_random.s1_xor_s0[18] ),
    .B(_04129_),
    .Y(_00009_));
 sky130_fd_sc_hd__xnor2_1 _09231_ (.A(\u_glbl_reg.u_random.s0[2] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[28] ),
    .Y(_04130_));
 sky130_fd_sc_hd__xnor2_1 _09232_ (.A(\u_glbl_reg.u_random.s1_xor_s0[19] ),
    .B(_04130_),
    .Y(_00010_));
 sky130_fd_sc_hd__xnor2_1 _09233_ (.A(\u_glbl_reg.u_random.s0[3] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[29] ),
    .Y(_04131_));
 sky130_fd_sc_hd__xnor2_1 _09234_ (.A(\u_glbl_reg.u_random.s1_xor_s0[20] ),
    .B(_04131_),
    .Y(_00012_));
 sky130_fd_sc_hd__xnor2_1 _09235_ (.A(\u_glbl_reg.u_random.s0[4] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[30] ),
    .Y(_04132_));
 sky130_fd_sc_hd__xnor2_1 _09236_ (.A(\u_glbl_reg.u_random.s1_xor_s0[21] ),
    .B(_04132_),
    .Y(_00013_));
 sky130_fd_sc_hd__xnor2_1 _09237_ (.A(\u_glbl_reg.u_random.s0[5] ),
    .B(\u_glbl_reg.u_random.s1_xor_s0[31] ),
    .Y(_04133_));
 sky130_fd_sc_hd__xnor2_1 _09238_ (.A(\u_glbl_reg.u_random.s1_xor_s0[22] ),
    .B(_04133_),
    .Y(_00014_));
 sky130_fd_sc_hd__o21ai_1 _09239_ (.A1(\u_glbl_reg.u_usb_clk_sel.A1 ),
    .A2(_01156_),
    .B1(_00244_),
    .Y(_00242_));
 sky130_fd_sc_hd__and2_1 _09240_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[0] ),
    .X(net333));
 sky130_fd_sc_hd__and2_1 _09241_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[1] ),
    .X(net344));
 sky130_fd_sc_hd__and2_1 _09242_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[2] ),
    .X(net355));
 sky130_fd_sc_hd__and2_1 _09243_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[3] ),
    .X(net358));
 sky130_fd_sc_hd__and2_1 _09244_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[4] ),
    .X(net359));
 sky130_fd_sc_hd__and2_1 _09245_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[5] ),
    .X(net360));
 sky130_fd_sc_hd__and2_1 _09246_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[6] ),
    .X(net361));
 sky130_fd_sc_hd__and2_1 _09247_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[7] ),
    .X(net362));
 sky130_fd_sc_hd__and2_2 _09248_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[8] ),
    .X(net363));
 sky130_fd_sc_hd__and2_1 _09249_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[9] ),
    .X(net364));
 sky130_fd_sc_hd__and2_1 _09250_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[10] ),
    .X(net334));
 sky130_fd_sc_hd__and2_1 _09251_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[11] ),
    .X(net335));
 sky130_fd_sc_hd__and2_1 _09252_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[12] ),
    .X(net336));
 sky130_fd_sc_hd__and2_1 _09253_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[13] ),
    .X(net337));
 sky130_fd_sc_hd__and2_1 _09254_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[14] ),
    .X(net338));
 sky130_fd_sc_hd__and2_1 _09255_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[15] ),
    .X(net339));
 sky130_fd_sc_hd__and2_1 _09256_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[16] ),
    .X(net340));
 sky130_fd_sc_hd__and2_2 _09257_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[17] ),
    .X(net341));
 sky130_fd_sc_hd__and2_2 _09258_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[18] ),
    .X(net342));
 sky130_fd_sc_hd__and2_2 _09259_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[19] ),
    .X(net343));
 sky130_fd_sc_hd__and2_2 _09260_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[20] ),
    .X(net345));
 sky130_fd_sc_hd__and2_2 _09261_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[21] ),
    .X(net346));
 sky130_fd_sc_hd__and2_1 _09262_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[22] ),
    .X(net347));
 sky130_fd_sc_hd__and2_1 _09263_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[23] ),
    .X(net348));
 sky130_fd_sc_hd__and2_1 _09264_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[24] ),
    .X(net349));
 sky130_fd_sc_hd__and2_1 _09265_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[25] ),
    .X(net350));
 sky130_fd_sc_hd__and2_1 _09266_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[26] ),
    .X(net351));
 sky130_fd_sc_hd__and2_1 _09267_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[27] ),
    .X(net352));
 sky130_fd_sc_hd__and2_1 _09268_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[28] ),
    .X(net353));
 sky130_fd_sc_hd__and2_1 _09269_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[29] ),
    .X(net354));
 sky130_fd_sc_hd__and2_1 _09270_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[30] ),
    .X(net356));
 sky130_fd_sc_hd__and2_1 _09271_ (.A(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ),
    .B(\u_glbl_reg.reg_3[31] ),
    .X(net357));
 sky130_fd_sc_hd__nand2_1 _09272_ (.A(\u_glbl_reg.u_random.n0[0] ),
    .B(\u_glbl_reg.u_random.n1[0] ),
    .Y(_04134_));
 sky130_fd_sc_hd__or2_1 _09273_ (.A(\u_glbl_reg.u_random.n0[0] ),
    .B(\u_glbl_reg.u_random.n1[0] ),
    .X(_04135_));
 sky130_fd_sc_hd__and2_1 _09274_ (.A(_04134_),
    .B(_04135_),
    .X(_00702_));
 sky130_fd_sc_hd__nand2_1 _09275_ (.A(\u_glbl_reg.u_random.n0[1] ),
    .B(\u_glbl_reg.u_random.n1[1] ),
    .Y(_04136_));
 sky130_fd_sc_hd__nor2_1 _09276_ (.A(\u_glbl_reg.u_random.n0[1] ),
    .B(\u_glbl_reg.u_random.n1[1] ),
    .Y(_04137_));
 sky130_fd_sc_hd__or2_1 _09277_ (.A(\u_glbl_reg.u_random.n0[1] ),
    .B(\u_glbl_reg.u_random.n1[1] ),
    .X(_04138_));
 sky130_fd_sc_hd__nand2_1 _09278_ (.A(_04136_),
    .B(_04138_),
    .Y(_04139_));
 sky130_fd_sc_hd__xor2_1 _09279_ (.A(_04134_),
    .B(_04139_),
    .X(_00713_));
 sky130_fd_sc_hd__o21a_1 _09280_ (.A1(_04134_),
    .A2(_04137_),
    .B1(_04136_),
    .X(_04140_));
 sky130_fd_sc_hd__nor2_1 _09281_ (.A(\u_glbl_reg.u_random.n0[2] ),
    .B(\u_glbl_reg.u_random.n1[2] ),
    .Y(_04141_));
 sky130_fd_sc_hd__nand2_1 _09282_ (.A(\u_glbl_reg.u_random.n0[2] ),
    .B(\u_glbl_reg.u_random.n1[2] ),
    .Y(_04142_));
 sky130_fd_sc_hd__and2b_1 _09283_ (.A_N(_04141_),
    .B(_04142_),
    .X(_04143_));
 sky130_fd_sc_hd__xnor2_1 _09284_ (.A(_04140_),
    .B(_04143_),
    .Y(_00724_));
 sky130_fd_sc_hd__nor2_1 _09285_ (.A(\u_glbl_reg.u_random.n0[3] ),
    .B(\u_glbl_reg.u_random.n1[3] ),
    .Y(_04144_));
 sky130_fd_sc_hd__nand2_1 _09286_ (.A(\u_glbl_reg.u_random.n0[3] ),
    .B(\u_glbl_reg.u_random.n1[3] ),
    .Y(_04145_));
 sky130_fd_sc_hd__nand2b_1 _09287_ (.A_N(_04144_),
    .B(_04145_),
    .Y(_04146_));
 sky130_fd_sc_hd__o21ai_1 _09288_ (.A1(_04140_),
    .A2(_04141_),
    .B1(_04142_),
    .Y(_04147_));
 sky130_fd_sc_hd__xnor2_1 _09289_ (.A(_04146_),
    .B(_04147_),
    .Y(_00727_));
 sky130_fd_sc_hd__or2_1 _09290_ (.A(\u_glbl_reg.u_random.n0[4] ),
    .B(\u_glbl_reg.u_random.n1[4] ),
    .X(_04148_));
 sky130_fd_sc_hd__nand2_1 _09291_ (.A(\u_glbl_reg.u_random.n0[4] ),
    .B(\u_glbl_reg.u_random.n1[4] ),
    .Y(_04149_));
 sky130_fd_sc_hd__nand2_1 _09292_ (.A(_04148_),
    .B(_04149_),
    .Y(_04150_));
 sky130_fd_sc_hd__o211a_1 _09293_ (.A1(_04140_),
    .A2(_04141_),
    .B1(_04142_),
    .C1(_04145_),
    .X(_04151_));
 sky130_fd_sc_hd__nor2_1 _09294_ (.A(_04144_),
    .B(_04151_),
    .Y(_04152_));
 sky130_fd_sc_hd__xnor2_1 _09295_ (.A(_04150_),
    .B(_04152_),
    .Y(_00728_));
 sky130_fd_sc_hd__or2_1 _09296_ (.A(\u_glbl_reg.u_random.n0[5] ),
    .B(\u_glbl_reg.u_random.n1[5] ),
    .X(_04153_));
 sky130_fd_sc_hd__nand2_1 _09297_ (.A(\u_glbl_reg.u_random.n0[5] ),
    .B(\u_glbl_reg.u_random.n1[5] ),
    .Y(_04154_));
 sky130_fd_sc_hd__nand2_1 _09298_ (.A(_04153_),
    .B(_04154_),
    .Y(_04155_));
 sky130_fd_sc_hd__o31ai_2 _09299_ (.A1(_04144_),
    .A2(_04150_),
    .A3(_04151_),
    .B1(_04149_),
    .Y(_04156_));
 sky130_fd_sc_hd__xnor2_1 _09300_ (.A(_04155_),
    .B(_04156_),
    .Y(_00729_));
 sky130_fd_sc_hd__or2_1 _09301_ (.A(\u_glbl_reg.u_random.n0[6] ),
    .B(\u_glbl_reg.u_random.n1[6] ),
    .X(_04157_));
 sky130_fd_sc_hd__nand2_1 _09302_ (.A(\u_glbl_reg.u_random.n0[6] ),
    .B(\u_glbl_reg.u_random.n1[6] ),
    .Y(_04158_));
 sky130_fd_sc_hd__nand2_1 _09303_ (.A(_04157_),
    .B(_04158_),
    .Y(_04159_));
 sky130_fd_sc_hd__a21boi_1 _09304_ (.A1(_04153_),
    .A2(_04156_),
    .B1_N(_04154_),
    .Y(_04160_));
 sky130_fd_sc_hd__xor2_1 _09305_ (.A(_04159_),
    .B(_04160_),
    .X(_00730_));
 sky130_fd_sc_hd__xnor2_1 _09306_ (.A(\u_glbl_reg.u_random.n0[7] ),
    .B(\u_glbl_reg.u_random.n1[7] ),
    .Y(_04161_));
 sky130_fd_sc_hd__o21ai_1 _09307_ (.A1(_04159_),
    .A2(_04160_),
    .B1(_04158_),
    .Y(_04162_));
 sky130_fd_sc_hd__xnor2_1 _09308_ (.A(_04161_),
    .B(_04162_),
    .Y(_00731_));
 sky130_fd_sc_hd__or2_1 _09309_ (.A(\u_glbl_reg.u_random.n0[8] ),
    .B(\u_glbl_reg.u_random.n1[8] ),
    .X(_04163_));
 sky130_fd_sc_hd__nand2_1 _09310_ (.A(\u_glbl_reg.u_random.n0[8] ),
    .B(\u_glbl_reg.u_random.n1[8] ),
    .Y(_04164_));
 sky130_fd_sc_hd__nand2_1 _09311_ (.A(_04163_),
    .B(_04164_),
    .Y(_04165_));
 sky130_fd_sc_hd__o211a_1 _09312_ (.A1(\u_glbl_reg.u_random.n0[7] ),
    .A2(\u_glbl_reg.u_random.n1[7] ),
    .B1(\u_glbl_reg.u_random.n1[6] ),
    .C1(\u_glbl_reg.u_random.n0[6] ),
    .X(_04166_));
 sky130_fd_sc_hd__a21oi_1 _09313_ (.A1(\u_glbl_reg.u_random.n0[7] ),
    .A2(\u_glbl_reg.u_random.n1[7] ),
    .B1(_04166_),
    .Y(_04167_));
 sky130_fd_sc_hd__o31a_1 _09314_ (.A1(_04159_),
    .A2(_04160_),
    .A3(_04161_),
    .B1(_04167_),
    .X(_04168_));
 sky130_fd_sc_hd__xor2_1 _09315_ (.A(_04165_),
    .B(_04168_),
    .X(_00732_));
 sky130_fd_sc_hd__nand2_1 _09316_ (.A(\u_glbl_reg.u_random.n0[9] ),
    .B(\u_glbl_reg.u_random.n1[9] ),
    .Y(_04169_));
 sky130_fd_sc_hd__inv_2 _09317_ (.A(_04169_),
    .Y(_04170_));
 sky130_fd_sc_hd__nor2_1 _09318_ (.A(\u_glbl_reg.u_random.n0[9] ),
    .B(\u_glbl_reg.u_random.n1[9] ),
    .Y(_04171_));
 sky130_fd_sc_hd__nor2_1 _09319_ (.A(_04170_),
    .B(_04171_),
    .Y(_04172_));
 sky130_fd_sc_hd__o21a_1 _09320_ (.A1(_04165_),
    .A2(_04168_),
    .B1(_04164_),
    .X(_04173_));
 sky130_fd_sc_hd__xnor2_1 _09321_ (.A(_04172_),
    .B(_04173_),
    .Y(_00733_));
 sky130_fd_sc_hd__or2_1 _09322_ (.A(\u_glbl_reg.u_random.n0[10] ),
    .B(\u_glbl_reg.u_random.n1[10] ),
    .X(_04174_));
 sky130_fd_sc_hd__nand2_1 _09323_ (.A(\u_glbl_reg.u_random.n0[10] ),
    .B(\u_glbl_reg.u_random.n1[10] ),
    .Y(_04175_));
 sky130_fd_sc_hd__nand2_1 _09324_ (.A(_04174_),
    .B(_04175_),
    .Y(_04176_));
 sky130_fd_sc_hd__o21ai_1 _09325_ (.A1(_04171_),
    .A2(_04173_),
    .B1(_04169_),
    .Y(_04177_));
 sky130_fd_sc_hd__xnor2_1 _09326_ (.A(_04176_),
    .B(_04177_),
    .Y(_00703_));
 sky130_fd_sc_hd__or2_1 _09327_ (.A(\u_glbl_reg.u_random.n0[11] ),
    .B(\u_glbl_reg.u_random.n1[11] ),
    .X(_04178_));
 sky130_fd_sc_hd__nand2_1 _09328_ (.A(\u_glbl_reg.u_random.n0[11] ),
    .B(\u_glbl_reg.u_random.n1[11] ),
    .Y(_04179_));
 sky130_fd_sc_hd__nand2_1 _09329_ (.A(_04178_),
    .B(_04179_),
    .Y(_04180_));
 sky130_fd_sc_hd__a21bo_1 _09330_ (.A1(_04174_),
    .A2(_04177_),
    .B1_N(_04175_),
    .X(_04181_));
 sky130_fd_sc_hd__xnor2_1 _09331_ (.A(_04180_),
    .B(_04181_),
    .Y(_00704_));
 sky130_fd_sc_hd__or2_1 _09332_ (.A(\u_glbl_reg.u_random.n0[12] ),
    .B(\u_glbl_reg.u_random.n1[12] ),
    .X(_04182_));
 sky130_fd_sc_hd__nand2_1 _09333_ (.A(\u_glbl_reg.u_random.n0[12] ),
    .B(\u_glbl_reg.u_random.n1[12] ),
    .Y(_04183_));
 sky130_fd_sc_hd__nand2_1 _09334_ (.A(_04182_),
    .B(_04183_),
    .Y(_04184_));
 sky130_fd_sc_hd__a2111o_1 _09335_ (.A1(_04164_),
    .A2(_04169_),
    .B1(_04171_),
    .C1(_04176_),
    .D1(_04180_),
    .X(_04185_));
 sky130_fd_sc_hd__nand2b_1 _09336_ (.A_N(_04175_),
    .B(_04178_),
    .Y(_04186_));
 sky130_fd_sc_hd__and3_1 _09337_ (.A(_04179_),
    .B(_04185_),
    .C(_04186_),
    .X(_04187_));
 sky130_fd_sc_hd__or3_1 _09338_ (.A(_04165_),
    .B(_04170_),
    .C(_04171_),
    .X(_04188_));
 sky130_fd_sc_hd__or3_1 _09339_ (.A(_04176_),
    .B(_04180_),
    .C(_04188_),
    .X(_04189_));
 sky130_fd_sc_hd__o21a_1 _09340_ (.A1(_04168_),
    .A2(_04189_),
    .B1(_04187_),
    .X(_04190_));
 sky130_fd_sc_hd__xor2_1 _09341_ (.A(_04184_),
    .B(_04190_),
    .X(_00705_));
 sky130_fd_sc_hd__and2_1 _09342_ (.A(\u_glbl_reg.u_random.n0[13] ),
    .B(\u_glbl_reg.u_random.n1[13] ),
    .X(_04191_));
 sky130_fd_sc_hd__nand2_1 _09343_ (.A(\u_glbl_reg.u_random.n0[13] ),
    .B(\u_glbl_reg.u_random.n1[13] ),
    .Y(_04192_));
 sky130_fd_sc_hd__nor2_1 _09344_ (.A(\u_glbl_reg.u_random.n0[13] ),
    .B(\u_glbl_reg.u_random.n1[13] ),
    .Y(_04193_));
 sky130_fd_sc_hd__nor2_1 _09345_ (.A(_04191_),
    .B(_04193_),
    .Y(_04194_));
 sky130_fd_sc_hd__o21a_1 _09346_ (.A1(_04184_),
    .A2(_04190_),
    .B1(_04183_),
    .X(_04195_));
 sky130_fd_sc_hd__xnor2_1 _09347_ (.A(_04194_),
    .B(_04195_),
    .Y(_00706_));
 sky130_fd_sc_hd__or2_1 _09348_ (.A(\u_glbl_reg.u_random.n0[14] ),
    .B(\u_glbl_reg.u_random.n1[14] ),
    .X(_04196_));
 sky130_fd_sc_hd__nand2_1 _09349_ (.A(\u_glbl_reg.u_random.n0[14] ),
    .B(\u_glbl_reg.u_random.n1[14] ),
    .Y(_04197_));
 sky130_fd_sc_hd__nand2_1 _09350_ (.A(_04196_),
    .B(_04197_),
    .Y(_04198_));
 sky130_fd_sc_hd__a21oi_1 _09351_ (.A1(_04192_),
    .A2(_04195_),
    .B1(_04193_),
    .Y(_04199_));
 sky130_fd_sc_hd__xnor2_1 _09352_ (.A(_04198_),
    .B(_04199_),
    .Y(_00707_));
 sky130_fd_sc_hd__nor2_1 _09353_ (.A(\u_glbl_reg.u_random.n0[15] ),
    .B(\u_glbl_reg.u_random.n1[15] ),
    .Y(_04200_));
 sky130_fd_sc_hd__nand2_1 _09354_ (.A(\u_glbl_reg.u_random.n0[15] ),
    .B(\u_glbl_reg.u_random.n1[15] ),
    .Y(_04201_));
 sky130_fd_sc_hd__nand2b_1 _09355_ (.A_N(_04200_),
    .B(_04201_),
    .Y(_04202_));
 sky130_fd_sc_hd__a21bo_1 _09356_ (.A1(_04196_),
    .A2(_04199_),
    .B1_N(_04197_),
    .X(_04203_));
 sky130_fd_sc_hd__xnor2_1 _09357_ (.A(_04202_),
    .B(_04203_),
    .Y(_00708_));
 sky130_fd_sc_hd__or3_1 _09358_ (.A(_04184_),
    .B(_04191_),
    .C(_04193_),
    .X(_04204_));
 sky130_fd_sc_hd__a31o_1 _09359_ (.A1(_04179_),
    .A2(_04185_),
    .A3(_04186_),
    .B1(_04204_),
    .X(_04205_));
 sky130_fd_sc_hd__o21a_1 _09360_ (.A1(_04183_),
    .A2(_04193_),
    .B1(_04192_),
    .X(_04206_));
 sky130_fd_sc_hd__a21bo_1 _09361_ (.A1(_04205_),
    .A2(_04206_),
    .B1_N(_04196_),
    .X(_04207_));
 sky130_fd_sc_hd__a31o_1 _09362_ (.A1(_04197_),
    .A2(_04201_),
    .A3(_04207_),
    .B1(_04200_),
    .X(_04208_));
 sky130_fd_sc_hd__or3_1 _09363_ (.A(_04198_),
    .B(_04202_),
    .C(_04204_),
    .X(_04209_));
 sky130_fd_sc_hd__o31a_2 _09364_ (.A1(_04168_),
    .A2(_04189_),
    .A3(_04209_),
    .B1(_04208_),
    .X(_04210_));
 sky130_fd_sc_hd__or2_1 _09365_ (.A(\u_glbl_reg.u_random.n0[16] ),
    .B(\u_glbl_reg.u_random.n1[16] ),
    .X(_04211_));
 sky130_fd_sc_hd__nand2_1 _09366_ (.A(\u_glbl_reg.u_random.n0[16] ),
    .B(\u_glbl_reg.u_random.n1[16] ),
    .Y(_04212_));
 sky130_fd_sc_hd__nand2_1 _09367_ (.A(_04211_),
    .B(_04212_),
    .Y(_04213_));
 sky130_fd_sc_hd__xor2_1 _09368_ (.A(_04210_),
    .B(_04213_),
    .X(_00709_));
 sky130_fd_sc_hd__nand2_1 _09369_ (.A(\u_glbl_reg.u_random.n0[17] ),
    .B(\u_glbl_reg.u_random.n1[17] ),
    .Y(_04214_));
 sky130_fd_sc_hd__inv_2 _09370_ (.A(_04214_),
    .Y(_04215_));
 sky130_fd_sc_hd__nor2_1 _09371_ (.A(\u_glbl_reg.u_random.n0[17] ),
    .B(\u_glbl_reg.u_random.n1[17] ),
    .Y(_04216_));
 sky130_fd_sc_hd__nor2_1 _09372_ (.A(_04215_),
    .B(_04216_),
    .Y(_04217_));
 sky130_fd_sc_hd__o21a_1 _09373_ (.A1(_04210_),
    .A2(_04213_),
    .B1(_04212_),
    .X(_04218_));
 sky130_fd_sc_hd__xnor2_1 _09374_ (.A(_04217_),
    .B(_04218_),
    .Y(_00710_));
 sky130_fd_sc_hd__or2_1 _09375_ (.A(\u_glbl_reg.u_random.n0[18] ),
    .B(\u_glbl_reg.u_random.n1[18] ),
    .X(_04219_));
 sky130_fd_sc_hd__and2_1 _09376_ (.A(\u_glbl_reg.u_random.n0[18] ),
    .B(\u_glbl_reg.u_random.n1[18] ),
    .X(_04220_));
 sky130_fd_sc_hd__xnor2_1 _09377_ (.A(\u_glbl_reg.u_random.n0[18] ),
    .B(\u_glbl_reg.u_random.n1[18] ),
    .Y(_04221_));
 sky130_fd_sc_hd__o21ai_1 _09378_ (.A1(_04216_),
    .A2(_04218_),
    .B1(_04214_),
    .Y(_04222_));
 sky130_fd_sc_hd__xnor2_1 _09379_ (.A(_04221_),
    .B(_04222_),
    .Y(_00711_));
 sky130_fd_sc_hd__xnor2_1 _09380_ (.A(\u_glbl_reg.u_random.n0[19] ),
    .B(\u_glbl_reg.u_random.n1[19] ),
    .Y(_04223_));
 sky130_fd_sc_hd__a21o_1 _09381_ (.A1(_04219_),
    .A2(_04222_),
    .B1(_04220_),
    .X(_04224_));
 sky130_fd_sc_hd__xnor2_1 _09382_ (.A(_04223_),
    .B(_04224_),
    .Y(_00712_));
 sky130_fd_sc_hd__or2_1 _09383_ (.A(\u_glbl_reg.u_random.n0[20] ),
    .B(\u_glbl_reg.u_random.n1[20] ),
    .X(_04225_));
 sky130_fd_sc_hd__nand2_1 _09384_ (.A(\u_glbl_reg.u_random.n0[20] ),
    .B(\u_glbl_reg.u_random.n1[20] ),
    .Y(_04226_));
 sky130_fd_sc_hd__nand2_1 _09385_ (.A(_04225_),
    .B(_04226_),
    .Y(_04227_));
 sky130_fd_sc_hd__or2_1 _09386_ (.A(_04221_),
    .B(_04223_),
    .X(_04228_));
 sky130_fd_sc_hd__a211oi_1 _09387_ (.A1(_04212_),
    .A2(_04214_),
    .B1(_04216_),
    .C1(_04228_),
    .Y(_04229_));
 sky130_fd_sc_hd__o21a_1 _09388_ (.A1(\u_glbl_reg.u_random.n0[19] ),
    .A2(\u_glbl_reg.u_random.n1[19] ),
    .B1(_04220_),
    .X(_04230_));
 sky130_fd_sc_hd__a211oi_1 _09389_ (.A1(\u_glbl_reg.u_random.n0[19] ),
    .A2(\u_glbl_reg.u_random.n1[19] ),
    .B1(_04229_),
    .C1(_04230_),
    .Y(_04231_));
 sky130_fd_sc_hd__or4_1 _09390_ (.A(_04213_),
    .B(_04215_),
    .C(_04216_),
    .D(_04228_),
    .X(_04232_));
 sky130_fd_sc_hd__o21ai_1 _09391_ (.A1(_04210_),
    .A2(_04232_),
    .B1(_04231_),
    .Y(_04233_));
 sky130_fd_sc_hd__xnor2_1 _09392_ (.A(_04227_),
    .B(_04233_),
    .Y(_00714_));
 sky130_fd_sc_hd__and2_1 _09393_ (.A(\u_glbl_reg.u_random.n0[21] ),
    .B(\u_glbl_reg.u_random.n1[21] ),
    .X(_04234_));
 sky130_fd_sc_hd__nand2_1 _09394_ (.A(\u_glbl_reg.u_random.n0[21] ),
    .B(\u_glbl_reg.u_random.n1[21] ),
    .Y(_04235_));
 sky130_fd_sc_hd__nor2_1 _09395_ (.A(\u_glbl_reg.u_random.n0[21] ),
    .B(\u_glbl_reg.u_random.n1[21] ),
    .Y(_04236_));
 sky130_fd_sc_hd__nor2_1 _09396_ (.A(_04234_),
    .B(_04236_),
    .Y(_04237_));
 sky130_fd_sc_hd__a21boi_1 _09397_ (.A1(_04225_),
    .A2(_04233_),
    .B1_N(_04226_),
    .Y(_04238_));
 sky130_fd_sc_hd__xnor2_1 _09398_ (.A(_04237_),
    .B(_04238_),
    .Y(_00715_));
 sky130_fd_sc_hd__nor2_1 _09399_ (.A(\u_glbl_reg.u_random.n0[22] ),
    .B(\u_glbl_reg.u_random.n1[22] ),
    .Y(_04239_));
 sky130_fd_sc_hd__nand2_1 _09400_ (.A(\u_glbl_reg.u_random.n0[22] ),
    .B(\u_glbl_reg.u_random.n1[22] ),
    .Y(_04240_));
 sky130_fd_sc_hd__nand2b_1 _09401_ (.A_N(_04239_),
    .B(_04240_),
    .Y(_04241_));
 sky130_fd_sc_hd__a21o_1 _09402_ (.A1(_04235_),
    .A2(_04238_),
    .B1(_04236_),
    .X(_04242_));
 sky130_fd_sc_hd__or2_1 _09403_ (.A(_04241_),
    .B(_04242_),
    .X(_04243_));
 sky130_fd_sc_hd__nand2_1 _09404_ (.A(_04241_),
    .B(_04242_),
    .Y(_04244_));
 sky130_fd_sc_hd__and2_1 _09405_ (.A(_04243_),
    .B(_04244_),
    .X(_00716_));
 sky130_fd_sc_hd__or2_1 _09406_ (.A(\u_glbl_reg.u_random.n0[23] ),
    .B(\u_glbl_reg.u_random.n1[23] ),
    .X(_04245_));
 sky130_fd_sc_hd__nand2_1 _09407_ (.A(\u_glbl_reg.u_random.n0[23] ),
    .B(\u_glbl_reg.u_random.n1[23] ),
    .Y(_04246_));
 sky130_fd_sc_hd__nand2_1 _09408_ (.A(_04245_),
    .B(_04246_),
    .Y(_04247_));
 sky130_fd_sc_hd__nand2_1 _09409_ (.A(_04240_),
    .B(_04243_),
    .Y(_04248_));
 sky130_fd_sc_hd__xnor2_1 _09410_ (.A(_04247_),
    .B(_04248_),
    .Y(_00717_));
 sky130_fd_sc_hd__or3_1 _09411_ (.A(_04227_),
    .B(_04234_),
    .C(_04236_),
    .X(_04249_));
 sky130_fd_sc_hd__o221a_1 _09412_ (.A1(_04226_),
    .A2(_04236_),
    .B1(_04249_),
    .B2(_04231_),
    .C1(_04235_),
    .X(_04250_));
 sky130_fd_sc_hd__o211ai_1 _09413_ (.A1(_04239_),
    .A2(_04250_),
    .B1(_04246_),
    .C1(_04240_),
    .Y(_04251_));
 sky130_fd_sc_hd__nand2_1 _09414_ (.A(_04245_),
    .B(_04251_),
    .Y(_04252_));
 sky130_fd_sc_hd__or3_1 _09415_ (.A(_04241_),
    .B(_04247_),
    .C(_04249_),
    .X(_04253_));
 sky130_fd_sc_hd__o31a_1 _09416_ (.A1(_04210_),
    .A2(_04232_),
    .A3(_04253_),
    .B1(_04252_),
    .X(_04254_));
 sky130_fd_sc_hd__nand2_1 _09417_ (.A(\u_glbl_reg.u_random.n0[24] ),
    .B(\u_glbl_reg.u_random.n1[24] ),
    .Y(_04255_));
 sky130_fd_sc_hd__or2_1 _09418_ (.A(\u_glbl_reg.u_random.n0[24] ),
    .B(\u_glbl_reg.u_random.n1[24] ),
    .X(_04256_));
 sky130_fd_sc_hd__nand2_1 _09419_ (.A(_04255_),
    .B(_04256_),
    .Y(_04257_));
 sky130_fd_sc_hd__xor2_1 _09420_ (.A(_04254_),
    .B(_04257_),
    .X(_00718_));
 sky130_fd_sc_hd__nand2_1 _09421_ (.A(\u_glbl_reg.u_random.n0[25] ),
    .B(\u_glbl_reg.u_random.n1[25] ),
    .Y(_04258_));
 sky130_fd_sc_hd__nor2_1 _09422_ (.A(\u_glbl_reg.u_random.n0[25] ),
    .B(\u_glbl_reg.u_random.n1[25] ),
    .Y(_04259_));
 sky130_fd_sc_hd__or2_1 _09423_ (.A(\u_glbl_reg.u_random.n0[25] ),
    .B(\u_glbl_reg.u_random.n1[25] ),
    .X(_04260_));
 sky130_fd_sc_hd__nand2_1 _09424_ (.A(_04258_),
    .B(_04260_),
    .Y(_04261_));
 sky130_fd_sc_hd__o21a_1 _09425_ (.A1(_04254_),
    .A2(_04257_),
    .B1(_04255_),
    .X(_04262_));
 sky130_fd_sc_hd__xor2_1 _09426_ (.A(_04261_),
    .B(_04262_),
    .X(_00719_));
 sky130_fd_sc_hd__or2_1 _09427_ (.A(\u_glbl_reg.u_random.n0[26] ),
    .B(\u_glbl_reg.u_random.n1[26] ),
    .X(_04263_));
 sky130_fd_sc_hd__nand2_1 _09428_ (.A(\u_glbl_reg.u_random.n0[26] ),
    .B(\u_glbl_reg.u_random.n1[26] ),
    .Y(_04264_));
 sky130_fd_sc_hd__nand2_1 _09429_ (.A(_04263_),
    .B(_04264_),
    .Y(_04265_));
 sky130_fd_sc_hd__a21oi_1 _09430_ (.A1(_04258_),
    .A2(_04262_),
    .B1(_04259_),
    .Y(_04266_));
 sky130_fd_sc_hd__xnor2_1 _09431_ (.A(_04265_),
    .B(_04266_),
    .Y(_00720_));
 sky130_fd_sc_hd__nor2_1 _09432_ (.A(\u_glbl_reg.u_random.n0[27] ),
    .B(\u_glbl_reg.u_random.n1[27] ),
    .Y(_04267_));
 sky130_fd_sc_hd__nand2_1 _09433_ (.A(\u_glbl_reg.u_random.n0[27] ),
    .B(\u_glbl_reg.u_random.n1[27] ),
    .Y(_04268_));
 sky130_fd_sc_hd__nand2b_1 _09434_ (.A_N(_04267_),
    .B(_04268_),
    .Y(_04269_));
 sky130_fd_sc_hd__a21bo_1 _09435_ (.A1(_04263_),
    .A2(_04266_),
    .B1_N(_04264_),
    .X(_04270_));
 sky130_fd_sc_hd__xnor2_1 _09436_ (.A(_04269_),
    .B(_04270_),
    .Y(_00721_));
 sky130_fd_sc_hd__or2_1 _09437_ (.A(_04265_),
    .B(_04269_),
    .X(_04271_));
 sky130_fd_sc_hd__or4_1 _09438_ (.A(_04254_),
    .B(_04257_),
    .C(_04261_),
    .D(_04271_),
    .X(_04272_));
 sky130_fd_sc_hd__a211o_1 _09439_ (.A1(_04255_),
    .A2(_04258_),
    .B1(_04259_),
    .C1(_04271_),
    .X(_04273_));
 sky130_fd_sc_hd__or2_1 _09440_ (.A(_04264_),
    .B(_04267_),
    .X(_04274_));
 sky130_fd_sc_hd__and4_1 _09441_ (.A(_04268_),
    .B(_04272_),
    .C(_04273_),
    .D(_04274_),
    .X(_04275_));
 sky130_fd_sc_hd__nor2_1 _09442_ (.A(\u_glbl_reg.u_random.n0[28] ),
    .B(\u_glbl_reg.u_random.n1[28] ),
    .Y(_04276_));
 sky130_fd_sc_hd__nand2_1 _09443_ (.A(\u_glbl_reg.u_random.n0[28] ),
    .B(\u_glbl_reg.u_random.n1[28] ),
    .Y(_04277_));
 sky130_fd_sc_hd__nand2b_1 _09444_ (.A_N(_04276_),
    .B(_04277_),
    .Y(_04278_));
 sky130_fd_sc_hd__xor2_1 _09445_ (.A(_04275_),
    .B(_04278_),
    .X(_00722_));
 sky130_fd_sc_hd__or2_1 _09446_ (.A(\u_glbl_reg.u_random.n0[29] ),
    .B(\u_glbl_reg.u_random.n1[29] ),
    .X(_04279_));
 sky130_fd_sc_hd__nand2_1 _09447_ (.A(\u_glbl_reg.u_random.n0[29] ),
    .B(\u_glbl_reg.u_random.n1[29] ),
    .Y(_04280_));
 sky130_fd_sc_hd__nand2_1 _09448_ (.A(_04279_),
    .B(_04280_),
    .Y(_04281_));
 sky130_fd_sc_hd__o21ai_1 _09449_ (.A1(_04275_),
    .A2(_04276_),
    .B1(_04277_),
    .Y(_04282_));
 sky130_fd_sc_hd__xnor2_1 _09450_ (.A(_04281_),
    .B(_04282_),
    .Y(_00723_));
 sky130_fd_sc_hd__nand2_1 _09451_ (.A(\u_glbl_reg.u_random.n0[30] ),
    .B(\u_glbl_reg.u_random.n1[30] ),
    .Y(_04283_));
 sky130_fd_sc_hd__or2_1 _09452_ (.A(\u_glbl_reg.u_random.n0[30] ),
    .B(\u_glbl_reg.u_random.n1[30] ),
    .X(_04284_));
 sky130_fd_sc_hd__nand2_1 _09453_ (.A(_04283_),
    .B(_04284_),
    .Y(_04285_));
 sky130_fd_sc_hd__a21bo_1 _09454_ (.A1(_04279_),
    .A2(_04282_),
    .B1_N(_04280_),
    .X(_04286_));
 sky130_fd_sc_hd__xnor2_1 _09455_ (.A(_04285_),
    .B(_04286_),
    .Y(_00725_));
 sky130_fd_sc_hd__a21bo_1 _09456_ (.A1(_04284_),
    .A2(_04286_),
    .B1_N(_04283_),
    .X(_04287_));
 sky130_fd_sc_hd__xnor2_2 _09457_ (.A(\u_glbl_reg.u_random.n0[31] ),
    .B(\u_glbl_reg.u_random.n1[31] ),
    .Y(_04288_));
 sky130_fd_sc_hd__xnor2_1 _09458_ (.A(_04287_),
    .B(_04288_),
    .Y(_00726_));
 sky130_fd_sc_hd__and2_1 _09459_ (.A(net1307),
    .B(net1374),
    .X(net384));
 sky130_fd_sc_hd__a31o_1 _09460_ (.A1(_00852_),
    .A2(net710),
    .A3(_01270_),
    .B1(_01559_),
    .X(_04289_));
 sky130_fd_sc_hd__a31o_1 _09461_ (.A1(_00850_),
    .A2(net714),
    .A3(_01270_),
    .B1(_00776_),
    .X(_04290_));
 sky130_fd_sc_hd__o21ba_1 _09462_ (.A1(_04289_),
    .A2(_04290_),
    .B1_N(_01560_),
    .X(_00578_));
 sky130_fd_sc_hd__and3_1 _09463_ (.A(net1337),
    .B(_01270_),
    .C(net1135),
    .X(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__nor2_1 _09464_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .B(_00849_),
    .Y(_00590_));
 sky130_fd_sc_hd__and2_1 _09465_ (.A(_04345_),
    .B(_00589_),
    .X(_00593_));
 sky130_fd_sc_hd__and2_1 _09466_ (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.wr_ptr ),
    .B(_00589_),
    .X(_00592_));
 sky130_fd_sc_hd__nor2_1 _09467_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ),
    .B(_00851_),
    .Y(_00583_));
 sky130_fd_sc_hd__and2_1 _09468_ (.A(_04343_),
    .B(_00582_),
    .X(_00586_));
 sky130_fd_sc_hd__and2_1 _09469_ (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.wr_ptr ),
    .B(_00582_),
    .X(_00585_));
 sky130_fd_sc_hd__and4_2 _09470_ (.A(net1335),
    .B(\u_pwm.reg_ack_glbl ),
    .C(net1158),
    .D(_01390_),
    .X(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ));
 sky130_fd_sc_hd__nand2_1 _09471_ (.A(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ),
    .B(_01040_),
    .Y(_04291_));
 sky130_fd_sc_hd__o21ba_1 _09472_ (.A1(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ),
    .A2(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .B1_N(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[2] ),
    .X(_04292_));
 sky130_fd_sc_hd__a32o_1 _09473_ (.A1(_00989_),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[2] ),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .B1(_04291_),
    .B2(_04292_),
    .X(_04293_));
 sky130_fd_sc_hd__mux4_1 _09474_ (.A0(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .A1(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .A2(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .S0(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ),
    .S1(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[2] ),
    .X(_04294_));
 sky130_fd_sc_hd__mux2_1 _09475_ (.A0(_04294_),
    .A1(_04293_),
    .S(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[1] ),
    .X(_04295_));
 sky130_fd_sc_hd__o21ai_1 _09476_ (.A1(\u_pwm.u_pwm_0.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_gpio_edge ),
    .B1(_04295_),
    .Y(_04296_));
 sky130_fd_sc_hd__a21o_1 _09477_ (.A1(\u_pwm.u_pwm_0.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_0.cfg_pwm_gpio_edge ),
    .B1(_04295_),
    .X(_04297_));
 sky130_fd_sc_hd__and4_1 _09478_ (.A(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_gpio_enb ),
    .C(_04296_),
    .D(_04297_),
    .X(_00318_));
 sky130_fd_sc_hd__and3_1 _09479_ (.A(\u_pwm.u_pwm_0.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_0.cfg_pwm_gpio_enb ),
    .C(_04295_),
    .X(_00317_));
 sky130_fd_sc_hd__nand2_1 _09480_ (.A(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ),
    .B(_01040_),
    .Y(_04298_));
 sky130_fd_sc_hd__o21ba_1 _09481_ (.A1(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ),
    .A2(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .B1_N(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[2] ),
    .X(_04299_));
 sky130_fd_sc_hd__a32o_1 _09482_ (.A1(_00990_),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[2] ),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .B1(_04298_),
    .B2(_04299_),
    .X(_04300_));
 sky130_fd_sc_hd__mux4_1 _09483_ (.A0(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .A1(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .A2(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .S0(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ),
    .S1(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[2] ),
    .X(_04301_));
 sky130_fd_sc_hd__mux2_1 _09484_ (.A0(_04301_),
    .A1(_04300_),
    .S(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[1] ),
    .X(_04302_));
 sky130_fd_sc_hd__o21ai_1 _09485_ (.A1(\u_pwm.u_pwm_1.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_gpio_edge ),
    .B1(_04302_),
    .Y(_04303_));
 sky130_fd_sc_hd__a21o_1 _09486_ (.A1(\u_pwm.u_pwm_1.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_1.cfg_pwm_gpio_edge ),
    .B1(_04302_),
    .X(_04304_));
 sky130_fd_sc_hd__and4_1 _09487_ (.A(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_gpio_enb ),
    .C(_04303_),
    .D(_04304_),
    .X(_00371_));
 sky130_fd_sc_hd__and3_1 _09488_ (.A(\u_pwm.u_pwm_1.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_1.cfg_pwm_gpio_enb ),
    .C(_04302_),
    .X(_00370_));
 sky130_fd_sc_hd__nand2_1 _09489_ (.A(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ),
    .B(_01040_),
    .Y(_04305_));
 sky130_fd_sc_hd__o21ba_1 _09490_ (.A1(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ),
    .A2(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .B1_N(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ),
    .X(_04306_));
 sky130_fd_sc_hd__a32o_1 _09491_ (.A1(_00991_),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ),
    .A3(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .B1(_04305_),
    .B2(_04306_),
    .X(_04307_));
 sky130_fd_sc_hd__mux4_2 _09492_ (.A0(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .A1(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .A2(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .A3(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .S0(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ),
    .S1(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ),
    .X(_04308_));
 sky130_fd_sc_hd__mux2_1 _09493_ (.A0(_04308_),
    .A1(_04307_),
    .S(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[1] ),
    .X(_04309_));
 sky130_fd_sc_hd__o21ai_1 _09494_ (.A1(\u_pwm.u_pwm_2.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_gpio_edge ),
    .B1(_04309_),
    .Y(_04310_));
 sky130_fd_sc_hd__a21o_1 _09495_ (.A1(\u_pwm.u_pwm_2.u_pwm.gpio_l ),
    .A2(\u_pwm.u_pwm_2.cfg_pwm_gpio_edge ),
    .B1(_04309_),
    .X(_04311_));
 sky130_fd_sc_hd__and4_1 _09496_ (.A(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_gpio_enb ),
    .C(_04310_),
    .D(_04311_),
    .X(_00424_));
 sky130_fd_sc_hd__and3_1 _09497_ (.A(\u_pwm.u_pwm_2.cfg_pwm_enb ),
    .B(\u_pwm.u_pwm_2.cfg_pwm_gpio_enb ),
    .C(_04309_),
    .X(_00423_));
 sky130_fd_sc_hd__nor2_1 _09498_ (.A(net1416),
    .B(_01561_),
    .Y(_04312_));
 sky130_fd_sc_hd__nand2_1 _09499_ (.A(net1300),
    .B(net1135),
    .Y(_04313_));
 sky130_fd_sc_hd__a2bb2o_1 _09500_ (.A1_N(\u_semaphore.reg_0[0] ),
    .A2_N(_04313_),
    .B1(net579),
    .B2(net1135),
    .X(_04314_));
 sky130_fd_sc_hd__a21o_1 _09501_ (.A1(\u_semaphore.reg_0[0] ),
    .A2(_04313_),
    .B1(_04314_),
    .X(_00734_));
 sky130_fd_sc_hd__nand2_1 _09502_ (.A(net1300),
    .B(net707),
    .Y(_04315_));
 sky130_fd_sc_hd__a2bb2o_1 _09503_ (.A1_N(\u_semaphore.reg_0[1] ),
    .A2_N(_04315_),
    .B1(net579),
    .B2(_01131_),
    .X(_04316_));
 sky130_fd_sc_hd__a21o_1 _09504_ (.A1(\u_semaphore.reg_0[1] ),
    .A2(_04315_),
    .B1(_04316_),
    .X(_00735_));
 sky130_fd_sc_hd__nand2_1 _09505_ (.A(net1300),
    .B(net697),
    .Y(_04317_));
 sky130_fd_sc_hd__a2bb2o_1 _09506_ (.A1_N(\u_semaphore.reg_0[2] ),
    .A2_N(_04317_),
    .B1(net579),
    .B2(net697),
    .X(_04318_));
 sky130_fd_sc_hd__a21o_1 _09507_ (.A1(\u_semaphore.reg_0[2] ),
    .A2(_04317_),
    .B1(_04318_),
    .X(_00736_));
 sky130_fd_sc_hd__nand2_1 _09508_ (.A(net1300),
    .B(net1140),
    .Y(_04319_));
 sky130_fd_sc_hd__a22oi_1 _09509_ (.A1(net1140),
    .A2(net579),
    .B1(_04319_),
    .B2(\u_semaphore.reg_0[3] ),
    .Y(_04320_));
 sky130_fd_sc_hd__o21ai_1 _09510_ (.A1(\u_semaphore.reg_0[3] ),
    .A2(_04319_),
    .B1(_04320_),
    .Y(_00737_));
 sky130_fd_sc_hd__and3_1 _09511_ (.A(net1300),
    .B(\u_semaphore.reg_0[4] ),
    .C(net711),
    .X(_04321_));
 sky130_fd_sc_hd__a21oi_1 _09512_ (.A1(net1301),
    .A2(net711),
    .B1(\u_semaphore.reg_0[4] ),
    .Y(_04322_));
 sky130_fd_sc_hd__a2bb2o_1 _09513_ (.A1_N(_04321_),
    .A2_N(_04322_),
    .B1(net711),
    .B2(net580),
    .X(_00738_));
 sky130_fd_sc_hd__nand2_1 _09514_ (.A(net1301),
    .B(_01001_),
    .Y(_04323_));
 sky130_fd_sc_hd__a22oi_1 _09515_ (.A1(_01001_),
    .A2(net580),
    .B1(_04323_),
    .B2(\u_semaphore.reg_0[5] ),
    .Y(_04324_));
 sky130_fd_sc_hd__o21ai_1 _09516_ (.A1(\u_semaphore.reg_0[5] ),
    .A2(_04323_),
    .B1(_04324_),
    .Y(_00739_));
 sky130_fd_sc_hd__nand2_1 _09517_ (.A(net1299),
    .B(net666),
    .Y(_04325_));
 sky130_fd_sc_hd__a2bb2o_1 _09518_ (.A1_N(\u_semaphore.reg_0[6] ),
    .A2_N(_04325_),
    .B1(net579),
    .B2(net667),
    .X(_04326_));
 sky130_fd_sc_hd__a21o_1 _09519_ (.A1(\u_semaphore.reg_0[6] ),
    .A2(_04325_),
    .B1(_04326_),
    .X(_00740_));
 sky130_fd_sc_hd__nand4_1 _09520_ (.A(net1300),
    .B(\u_semaphore.reg_0[7] ),
    .C(net1182),
    .D(net1145),
    .Y(_04327_));
 sky130_fd_sc_hd__a31o_1 _09521_ (.A1(net1300),
    .A2(net1182),
    .A3(net1145),
    .B1(\u_semaphore.reg_0[7] ),
    .X(_04328_));
 sky130_fd_sc_hd__a22o_1 _09522_ (.A1(net670),
    .A2(net579),
    .B1(_04327_),
    .B2(_04328_),
    .X(_00741_));
 sky130_fd_sc_hd__and2_1 _09523_ (.A(net1564),
    .B(net774),
    .X(_00742_));
 sky130_fd_sc_hd__and2_1 _09524_ (.A(net1556),
    .B(net774),
    .X(_00743_));
 sky130_fd_sc_hd__and2_1 _09525_ (.A(net1549),
    .B(net781),
    .X(_00744_));
 sky130_fd_sc_hd__and2_1 _09526_ (.A(net1541),
    .B(net774),
    .X(_00745_));
 sky130_fd_sc_hd__and2_1 _09527_ (.A(net1425),
    .B(net787),
    .X(_00746_));
 sky130_fd_sc_hd__and2_1 _09528_ (.A(net1418),
    .B(net780),
    .X(_00747_));
 sky130_fd_sc_hd__and2_1 _09529_ (.A(net1286),
    .B(net777),
    .X(_00748_));
 sky130_fd_sc_hd__and2_1 _09530_ (.A(net1645),
    .B(net782),
    .X(_00749_));
 sky130_fd_sc_hd__and2_1 _09531_ (.A(net1638),
    .B(net773),
    .X(_00750_));
 sky130_fd_sc_hd__and2_1 _09532_ (.A(net1628),
    .B(net785),
    .X(_00751_));
 sky130_fd_sc_hd__and2_1 _09533_ (.A(net1623),
    .B(net777),
    .X(_00752_));
 sky130_fd_sc_hd__and2_1 _09534_ (.A(net1614),
    .B(net787),
    .X(_00753_));
 sky130_fd_sc_hd__and2_1 _09535_ (.A(net1293),
    .B(net740),
    .X(_00754_));
 sky130_fd_sc_hd__and2_1 _09536_ (.A(net1572),
    .B(net752),
    .X(_00755_));
 sky130_fd_sc_hd__and2_1 _09537_ (.A(net1488),
    .B(net743),
    .X(_00756_));
 sky130_fd_sc_hd__and2_1 _09538_ (.A(net1466),
    .B(net742),
    .X(_00757_));
 sky130_fd_sc_hd__and2_1 _09539_ (.A(net1457),
    .B(net742),
    .X(_00758_));
 sky130_fd_sc_hd__and2_1 _09540_ (.A(net1448),
    .B(net740),
    .X(_00759_));
 sky130_fd_sc_hd__and2_1 _09541_ (.A(net1441),
    .B(net743),
    .X(_00760_));
 sky130_fd_sc_hd__and2_1 _09542_ (.A(net1433),
    .B(net752),
    .X(_00761_));
 sky130_fd_sc_hd__nand2_1 _09543_ (.A(net1299),
    .B(net662),
    .Y(_04329_));
 sky130_fd_sc_hd__a22oi_1 _09544_ (.A1(net662),
    .A2(net579),
    .B1(_04329_),
    .B2(\u_semaphore.reg_0[8] ),
    .Y(_04330_));
 sky130_fd_sc_hd__o21ai_1 _09545_ (.A1(\u_semaphore.reg_0[8] ),
    .A2(_04329_),
    .B1(_04330_),
    .Y(_00762_));
 sky130_fd_sc_hd__nand4_1 _09546_ (.A(net1299),
    .B(\u_semaphore.reg_0[9] ),
    .C(net1179),
    .D(net1152),
    .Y(_04331_));
 sky130_fd_sc_hd__a31o_1 _09547_ (.A1(net1299),
    .A2(net1179),
    .A3(net1152),
    .B1(\u_semaphore.reg_0[9] ),
    .X(_04332_));
 sky130_fd_sc_hd__a32o_1 _09548_ (.A1(net1179),
    .A2(net1152),
    .A3(net579),
    .B1(_04331_),
    .B2(_04332_),
    .X(_00763_));
 sky130_fd_sc_hd__nand4_1 _09549_ (.A(net1299),
    .B(\u_semaphore.reg_0[10] ),
    .C(net1160),
    .D(net1152),
    .Y(_04333_));
 sky130_fd_sc_hd__a31o_1 _09550_ (.A1(net1299),
    .A2(net1160),
    .A3(net1152),
    .B1(\u_semaphore.reg_0[10] ),
    .X(_04334_));
 sky130_fd_sc_hd__a32o_1 _09551_ (.A1(net1160),
    .A2(net1152),
    .A3(net579),
    .B1(_04333_),
    .B2(_04334_),
    .X(_00764_));
 sky130_fd_sc_hd__and3_1 _09552_ (.A(net1299),
    .B(net1152),
    .C(net1146),
    .X(_04335_));
 sky130_fd_sc_hd__xor2_1 _09553_ (.A(\u_semaphore.reg_0[11] ),
    .B(_04335_),
    .X(_04336_));
 sky130_fd_sc_hd__a31o_1 _09554_ (.A1(net1152),
    .A2(net1146),
    .A3(net579),
    .B1(_04336_),
    .X(_00765_));
 sky130_fd_sc_hd__and3_1 _09555_ (.A(net1299),
    .B(net1249),
    .C(_01144_),
    .X(_04337_));
 sky130_fd_sc_hd__xor2_1 _09556_ (.A(\u_semaphore.reg_0[12] ),
    .B(_04337_),
    .X(_04338_));
 sky130_fd_sc_hd__a31o_1 _09557_ (.A1(net1249),
    .A2(_01144_),
    .A3(net580),
    .B1(_04338_),
    .X(_00766_));
 sky130_fd_sc_hd__and3_1 _09558_ (.A(net1299),
    .B(net1180),
    .C(_01144_),
    .X(_04339_));
 sky130_fd_sc_hd__xor2_1 _09559_ (.A(\u_semaphore.reg_0[13] ),
    .B(_04339_),
    .X(_04340_));
 sky130_fd_sc_hd__a31o_1 _09560_ (.A1(net1180),
    .A2(_01144_),
    .A3(net580),
    .B1(_04340_),
    .X(_00767_));
 sky130_fd_sc_hd__and3_1 _09561_ (.A(net1301),
    .B(net1160),
    .C(_01144_),
    .X(_04341_));
 sky130_fd_sc_hd__xor2_1 _09562_ (.A(\u_semaphore.reg_0[14] ),
    .B(_04341_),
    .X(_04342_));
 sky130_fd_sc_hd__a31o_1 _09563_ (.A1(net1161),
    .A2(_01144_),
    .A3(net580),
    .B1(_04342_),
    .X(_00768_));
 sky130_fd_sc_hd__and2_1 _09564_ (.A(net1534),
    .B(net735),
    .X(_00770_));
 sky130_fd_sc_hd__and2_1 _09565_ (.A(net1526),
    .B(net735),
    .X(_00771_));
 sky130_fd_sc_hd__and2_1 _09566_ (.A(net1505),
    .B(net735),
    .X(_00772_));
 sky130_fd_sc_hd__and2_1 _09567_ (.A(net1498),
    .B(net735),
    .X(_00773_));
 sky130_fd_sc_hd__and2_1 _09568_ (.A(net1481),
    .B(net735),
    .X(_00774_));
 sky130_fd_sc_hd__nor2_1 _09569_ (.A(_01179_),
    .B(_01196_),
    .Y(_00646_));
 sky130_fd_sc_hd__a21oi_1 _09570_ (.A1(\u_ws281x.u_txd_1.state ),
    .A2(_01236_),
    .B1(_01221_),
    .Y(_00697_));
 sky130_fd_sc_hd__clkbuf_1 _09571_ (.A(\u_semaphore.reg_0[15] ),
    .X(_00769_));
 sky130_fd_sc_hd__dfrtp_1 _09572_ (.CLK(clknet_leaf_80_mclk),
    .D(net1346),
    .RESET_B(net976),
    .Q(\u_pwm.blk_sel[0] ));
 sky130_fd_sc_hd__dfrtp_4 _09573_ (.CLK(clknet_leaf_104_mclk),
    .D(net1345),
    .RESET_B(net857),
    .Q(\u_pwm.blk_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09574_ (.CLK(clknet_leaf_80_mclk),
    .D(net1344),
    .RESET_B(net976),
    .Q(\u_pwm.blk_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09575_ (.CLK(clknet_leaf_128_mclk),
    .D(net1689),
    .RESET_B(net48),
    .Q(\u_prst_sync.in_data_s ));
 sky130_fd_sc_hd__conb_1 _09575__1689 (.HI(net1689));
 sky130_fd_sc_hd__dfrtp_1 _09576_ (.CLK(clknet_leaf_128_mclk),
    .D(net2306),
    .RESET_B(net48),
    .Q(\u_prst_sync.in_data_2s ));
 sky130_fd_sc_hd__dfxtp_1 _09577_ (.CLK(clknet_1_1__leaf__04419_),
    .D(_00036_),
    .Q(\u_glbl_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfxtp_1 _09578_ (.CLK(clknet_1_1__leaf__04419_),
    .D(_00037_),
    .Q(\u_glbl_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09579_ (.CLK(clknet_1_0__leaf__04630_),
    .D(_00734_),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09580_ (.CLK(clknet_1_0__leaf__04630_),
    .D(_00735_),
    .RESET_B(net989),
    .Q(\u_semaphore.reg_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09581_ (.CLK(clknet_1_1__leaf__04630_),
    .D(_00736_),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09582_ (.CLK(clknet_1_1__leaf__04630_),
    .D(_00737_),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09583_ (.CLK(clknet_1_1__leaf__04630_),
    .D(_00738_),
    .RESET_B(net989),
    .Q(\u_semaphore.reg_0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _09584_ (.CLK(clknet_1_1__leaf__04630_),
    .D(_00739_),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_0[5] ));
 sky130_fd_sc_hd__dfrtp_2 _09585_ (.CLK(clknet_1_0__leaf__04630_),
    .D(_00740_),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09586_ (.CLK(clknet_1_0__leaf__04630_),
    .D(_00741_),
    .RESET_B(net988),
    .Q(\u_semaphore.reg_0[7] ));
 sky130_fd_sc_hd__dfxtp_2 _09587_ (.CLK(clknet_1_0__leaf__04418_),
    .D(_00032_),
    .Q(\u_glbl_reg.reg_2[16] ));
 sky130_fd_sc_hd__dfxtp_2 _09588_ (.CLK(clknet_1_0__leaf__04418_),
    .D(_00033_),
    .Q(\u_glbl_reg.reg_2[17] ));
 sky130_fd_sc_hd__dfxtp_4 _09589_ (.CLK(clknet_1_0__leaf__04418_),
    .D(_00034_),
    .Q(\u_glbl_reg.reg_2[18] ));
 sky130_fd_sc_hd__dfxtp_2 _09590_ (.CLK(clknet_1_0__leaf__04418_),
    .D(_00035_),
    .Q(\u_glbl_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_2 _09591_ (.CLK(clknet_leaf_81_mclk),
    .D(\u_gpio.u_bit[0].u_dglitch.gpio_out ),
    .RESET_B(net877),
    .Q(\u_gpio.u_bit[0].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09592_ (.CLK(clknet_leaf_104_mclk),
    .D(\u_gpio.u_bit[1].u_dglitch.gpio_out ),
    .RESET_B(net857),
    .Q(\u_gpio.u_bit[1].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09593_ (.CLK(clknet_leaf_81_mclk),
    .D(\u_gpio.u_bit[2].u_dglitch.gpio_out ),
    .RESET_B(net875),
    .Q(\u_gpio.u_bit[2].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09594_ (.CLK(clknet_leaf_106_mclk),
    .D(\u_gpio.u_bit[3].u_dglitch.gpio_out ),
    .RESET_B(net809),
    .Q(\u_gpio.u_bit[3].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_2 _09595_ (.CLK(clknet_leaf_90_mclk),
    .D(\u_gpio.u_bit[4].u_dglitch.gpio_out ),
    .RESET_B(net892),
    .Q(\u_gpio.u_bit[4].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09596_ (.CLK(clknet_leaf_16_mclk),
    .D(\u_gpio.u_bit[8].u_dglitch.gpio_out ),
    .RESET_B(net811),
    .Q(\u_gpio.u_bit[8].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09597_ (.CLK(clknet_leaf_107_mclk),
    .D(\u_gpio.u_bit[9].u_dglitch.gpio_out ),
    .RESET_B(net798),
    .Q(\u_gpio.u_bit[9].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09598_ (.CLK(clknet_leaf_110_mclk),
    .D(\u_gpio.u_bit[10].u_dglitch.gpio_out ),
    .RESET_B(net793),
    .Q(\u_gpio.u_bit[10].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09599_ (.CLK(clknet_leaf_11_mclk),
    .D(\u_gpio.u_bit[11].u_dglitch.gpio_out ),
    .RESET_B(net792),
    .Q(\u_gpio.u_bit[11].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09600_ (.CLK(clknet_leaf_15_mclk),
    .D(\u_gpio.u_bit[12].u_dglitch.gpio_out ),
    .RESET_B(net810),
    .Q(\u_gpio.u_bit[12].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09601_ (.CLK(clknet_leaf_13_mclk),
    .D(\u_gpio.u_bit[13].u_dglitch.gpio_out ),
    .RESET_B(net803),
    .Q(\u_gpio.u_bit[13].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09602_ (.CLK(clknet_leaf_14_mclk),
    .D(\u_gpio.u_bit[14].u_dglitch.gpio_out ),
    .RESET_B(net804),
    .Q(\u_gpio.u_bit[14].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09603_ (.CLK(clknet_leaf_19_mclk),
    .D(\u_gpio.u_bit[15].u_dglitch.gpio_out ),
    .RESET_B(net916),
    .Q(\u_gpio.u_bit[15].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_4 _09604_ (.CLK(clknet_leaf_17_mclk),
    .D(\u_gpio.u_bit[16].u_dglitch.gpio_out ),
    .RESET_B(net923),
    .Q(\u_gpio.u_bit[16].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_4 _09605_ (.CLK(clknet_leaf_79_mclk),
    .D(\u_gpio.u_bit[17].u_dglitch.gpio_out ),
    .RESET_B(net979),
    .Q(\u_gpio.u_bit[17].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09606_ (.CLK(clknet_leaf_20_mclk),
    .D(\u_gpio.u_bit[18].u_dglitch.gpio_out ),
    .RESET_B(net917),
    .Q(\u_gpio.u_bit[18].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09607_ (.CLK(clknet_leaf_22_mclk),
    .D(\u_gpio.u_bit[19].u_dglitch.gpio_out ),
    .RESET_B(net926),
    .Q(\u_gpio.u_bit[19].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_2 _09608_ (.CLK(clknet_leaf_53_mclk),
    .D(\u_gpio.u_bit[20].u_dglitch.gpio_out ),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[20].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09609_ (.CLK(clknet_leaf_22_mclk),
    .D(\u_gpio.u_bit[21].u_dglitch.gpio_out ),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[21].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09610_ (.CLK(clknet_leaf_17_mclk),
    .D(\u_gpio.u_bit[22].u_dglitch.gpio_out ),
    .RESET_B(net921),
    .Q(\u_gpio.u_bit[22].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_2 _09611_ (.CLK(clknet_leaf_115_mclk),
    .D(\u_gpio.u_bit[24].u_dglitch.gpio_out ),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[24].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_4 _09612_ (.CLK(clknet_leaf_92_mclk),
    .D(\u_gpio.u_bit[25].u_dglitch.gpio_out ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[25].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09613_ (.CLK(clknet_leaf_114_mclk),
    .D(\u_gpio.u_bit[26].u_dglitch.gpio_out ),
    .RESET_B(net767),
    .Q(\u_gpio.u_bit[26].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_4 _09614_ (.CLK(clknet_leaf_92_mclk),
    .D(\u_gpio.u_bit[27].u_dglitch.gpio_out ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[27].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_4 _09615_ (.CLK(clknet_leaf_103_mclk),
    .D(\u_gpio.u_bit[28].u_dglitch.gpio_out ),
    .RESET_B(net852),
    .Q(\u_gpio.u_bit[28].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09616_ (.CLK(clknet_leaf_112_mclk),
    .D(\u_gpio.u_bit[29].u_dglitch.gpio_out ),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[29].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09617_ (.CLK(clknet_leaf_112_mclk),
    .D(\u_gpio.u_bit[30].u_dglitch.gpio_out ),
    .RESET_B(net768),
    .Q(\u_gpio.u_bit[30].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_2 _09618_ (.CLK(clknet_leaf_115_mclk),
    .D(\u_gpio.u_bit[31].u_dglitch.gpio_out ),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[31].u_dglitch.gpio_reg ));
 sky130_fd_sc_hd__dfrtp_1 _09619_ (.CLK(clknet_1_0__leaf__04465_),
    .D(net1392),
    .RESET_B(net893),
    .Q(\u_gpio.u_bit[0].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09620_ (.CLK(clknet_1_1__leaf__04465_),
    .D(net2246),
    .RESET_B(net894),
    .Q(\u_gpio.u_bit[0].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09621_ (.CLK(clknet_1_1__leaf__04465_),
    .D(\u_gpio.u_bit[0].u_dglitch.gpio_ss[1] ),
    .RESET_B(net893),
    .Q(\u_gpio.u_bit[0].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09622_ (.CLK(clknet_1_0__leaf__04465_),
    .D(\u_gpio.u_bit[0].u_dglitch.gpio_ss[2] ),
    .RESET_B(net893),
    .Q(\u_gpio.u_bit[0].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09623_ (.CLK(clknet_1_1__leaf__04466_),
    .D(net1497),
    .RESET_B(net791),
    .Q(\u_gpio.u_bit[10].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09624_ (.CLK(clknet_1_0__leaf__04466_),
    .D(net2257),
    .RESET_B(net791),
    .Q(\u_gpio.u_bit[10].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09625_ (.CLK(clknet_1_1__leaf__04466_),
    .D(\u_gpio.u_bit[10].u_dglitch.gpio_ss[1] ),
    .RESET_B(net791),
    .Q(\u_gpio.u_bit[10].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09626_ (.CLK(clknet_1_0__leaf__04466_),
    .D(\u_gpio.u_bit[10].u_dglitch.gpio_ss[2] ),
    .RESET_B(net791),
    .Q(\u_gpio.u_bit[10].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09627_ (.CLK(clknet_1_1__leaf__04467_),
    .D(net1417),
    .RESET_B(net792),
    .Q(\u_gpio.u_bit[11].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09628_ (.CLK(clknet_1_1__leaf__04467_),
    .D(net2305),
    .RESET_B(net792),
    .Q(\u_gpio.u_bit[11].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09629_ (.CLK(clknet_1_0__leaf__04467_),
    .D(\u_gpio.u_bit[11].u_dglitch.gpio_ss[1] ),
    .RESET_B(net792),
    .Q(\u_gpio.u_bit[11].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09630_ (.CLK(clknet_1_0__leaf__04467_),
    .D(\u_gpio.u_bit[11].u_dglitch.gpio_ss[2] ),
    .RESET_B(net792),
    .Q(\u_gpio.u_bit[11].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09631_ (.CLK(clknet_1_0__leaf__04468_),
    .D(net1403),
    .RESET_B(net808),
    .Q(\u_gpio.u_bit[12].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09632_ (.CLK(clknet_1_1__leaf__04468_),
    .D(net2265),
    .RESET_B(net808),
    .Q(\u_gpio.u_bit[12].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09633_ (.CLK(clknet_1_1__leaf__04468_),
    .D(\u_gpio.u_bit[12].u_dglitch.gpio_ss[1] ),
    .RESET_B(net808),
    .Q(\u_gpio.u_bit[12].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09634_ (.CLK(clknet_1_0__leaf__04468_),
    .D(\u_gpio.u_bit[12].u_dglitch.gpio_ss[2] ),
    .RESET_B(net808),
    .Q(\u_gpio.u_bit[12].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09635_ (.CLK(clknet_1_0__leaf__04469_),
    .D(net1400),
    .RESET_B(net803),
    .Q(\u_gpio.u_bit[13].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09636_ (.CLK(clknet_1_0__leaf__04469_),
    .D(net2285),
    .RESET_B(net803),
    .Q(\u_gpio.u_bit[13].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09637_ (.CLK(clknet_1_1__leaf__04469_),
    .D(\u_gpio.u_bit[13].u_dglitch.gpio_ss[1] ),
    .RESET_B(net801),
    .Q(\u_gpio.u_bit[13].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09638_ (.CLK(clknet_1_1__leaf__04469_),
    .D(\u_gpio.u_bit[13].u_dglitch.gpio_ss[2] ),
    .RESET_B(net801),
    .Q(\u_gpio.u_bit[13].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09639_ (.CLK(clknet_1_0__leaf__04470_),
    .D(net1375),
    .RESET_B(net787),
    .Q(\u_gpio.u_bit[14].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09640_ (.CLK(clknet_1_1__leaf__04470_),
    .D(net2260),
    .RESET_B(net786),
    .Q(\u_gpio.u_bit[14].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09641_ (.CLK(clknet_1_1__leaf__04470_),
    .D(\u_gpio.u_bit[14].u_dglitch.gpio_ss[1] ),
    .RESET_B(net804),
    .Q(\u_gpio.u_bit[14].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09642_ (.CLK(clknet_1_0__leaf__04470_),
    .D(\u_gpio.u_bit[14].u_dglitch.gpio_ss[2] ),
    .RESET_B(net804),
    .Q(\u_gpio.u_bit[14].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09643_ (.CLK(clknet_1_0__leaf__04471_),
    .D(net1339),
    .RESET_B(net916),
    .Q(\u_gpio.u_bit[15].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09644_ (.CLK(clknet_1_1__leaf__04471_),
    .D(net2264),
    .RESET_B(net916),
    .Q(\u_gpio.u_bit[15].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09645_ (.CLK(clknet_1_0__leaf__04471_),
    .D(\u_gpio.u_bit[15].u_dglitch.gpio_ss[1] ),
    .RESET_B(net916),
    .Q(\u_gpio.u_bit[15].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09646_ (.CLK(clknet_1_1__leaf__04471_),
    .D(\u_gpio.u_bit[15].u_dglitch.gpio_ss[2] ),
    .RESET_B(net916),
    .Q(\u_gpio.u_bit[15].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09647_ (.CLK(clknet_1_0__leaf__04472_),
    .D(net17),
    .RESET_B(net1011),
    .Q(\u_gpio.u_bit[16].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09648_ (.CLK(clknet_1_0__leaf__04472_),
    .D(net2273),
    .RESET_B(net1007),
    .Q(\u_gpio.u_bit[16].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09649_ (.CLK(clknet_1_1__leaf__04472_),
    .D(\u_gpio.u_bit[16].u_dglitch.gpio_ss[1] ),
    .RESET_B(net1007),
    .Q(\u_gpio.u_bit[16].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09650_ (.CLK(clknet_1_1__leaf__04472_),
    .D(\u_gpio.u_bit[16].u_dglitch.gpio_ss[2] ),
    .RESET_B(net1007),
    .Q(\u_gpio.u_bit[16].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09651_ (.CLK(clknet_1_1__leaf__04473_),
    .D(net18),
    .RESET_B(net1008),
    .Q(\u_gpio.u_bit[17].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09652_ (.CLK(clknet_1_1__leaf__04473_),
    .D(net2287),
    .RESET_B(net1008),
    .Q(\u_gpio.u_bit[17].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09653_ (.CLK(clknet_1_0__leaf__04473_),
    .D(\u_gpio.u_bit[17].u_dglitch.gpio_ss[1] ),
    .RESET_B(net1008),
    .Q(\u_gpio.u_bit[17].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09654_ (.CLK(clknet_1_0__leaf__04473_),
    .D(\u_gpio.u_bit[17].u_dglitch.gpio_ss[2] ),
    .RESET_B(net1008),
    .Q(\u_gpio.u_bit[17].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09655_ (.CLK(clknet_1_0__leaf__04474_),
    .D(net19),
    .RESET_B(net904),
    .Q(\u_gpio.u_bit[18].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09656_ (.CLK(clknet_1_0__leaf__04474_),
    .D(net2281),
    .RESET_B(net904),
    .Q(\u_gpio.u_bit[18].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09657_ (.CLK(clknet_1_1__leaf__04474_),
    .D(\u_gpio.u_bit[18].u_dglitch.gpio_ss[1] ),
    .RESET_B(net904),
    .Q(\u_gpio.u_bit[18].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09658_ (.CLK(clknet_1_1__leaf__04474_),
    .D(\u_gpio.u_bit[18].u_dglitch.gpio_ss[2] ),
    .RESET_B(net904),
    .Q(\u_gpio.u_bit[18].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09659_ (.CLK(clknet_1_0__leaf__04475_),
    .D(net20),
    .RESET_B(net911),
    .Q(\u_gpio.u_bit[19].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09660_ (.CLK(clknet_1_0__leaf__04475_),
    .D(net2283),
    .RESET_B(net910),
    .Q(\u_gpio.u_bit[19].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09661_ (.CLK(clknet_1_1__leaf__04475_),
    .D(\u_gpio.u_bit[19].u_dglitch.gpio_ss[1] ),
    .RESET_B(net911),
    .Q(\u_gpio.u_bit[19].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09662_ (.CLK(clknet_1_1__leaf__04475_),
    .D(\u_gpio.u_bit[19].u_dglitch.gpio_ss[2] ),
    .RESET_B(net910),
    .Q(\u_gpio.u_bit[19].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09663_ (.CLK(clknet_1_1__leaf__04476_),
    .D(net14),
    .RESET_B(net800),
    .Q(\u_gpio.u_bit[1].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09664_ (.CLK(clknet_1_0__leaf__04476_),
    .D(net2236),
    .RESET_B(net800),
    .Q(\u_gpio.u_bit[1].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09665_ (.CLK(clknet_1_0__leaf__04476_),
    .D(\u_gpio.u_bit[1].u_dglitch.gpio_ss[1] ),
    .RESET_B(net799),
    .Q(\u_gpio.u_bit[1].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09666_ (.CLK(clknet_1_1__leaf__04476_),
    .D(\u_gpio.u_bit[1].u_dglitch.gpio_ss[2] ),
    .RESET_B(net799),
    .Q(\u_gpio.u_bit[1].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09667_ (.CLK(clknet_1_0__leaf__04477_),
    .D(net21),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[20].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09668_ (.CLK(clknet_1_1__leaf__04477_),
    .D(net2252),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[20].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09669_ (.CLK(clknet_1_0__leaf__04477_),
    .D(\u_gpio.u_bit[20].u_dglitch.gpio_ss[1] ),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[20].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09670_ (.CLK(clknet_1_1__leaf__04477_),
    .D(\u_gpio.u_bit[20].u_dglitch.gpio_ss[2] ),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[20].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09671_ (.CLK(clknet_1_0__leaf__04478_),
    .D(net22),
    .RESET_B(net913),
    .Q(\u_gpio.u_bit[21].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09672_ (.CLK(clknet_1_0__leaf__04478_),
    .D(net2297),
    .RESET_B(net913),
    .Q(\u_gpio.u_bit[21].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09673_ (.CLK(clknet_1_1__leaf__04478_),
    .D(\u_gpio.u_bit[21].u_dglitch.gpio_ss[1] ),
    .RESET_B(net913),
    .Q(\u_gpio.u_bit[21].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09674_ (.CLK(clknet_1_1__leaf__04478_),
    .D(\u_gpio.u_bit[21].u_dglitch.gpio_ss[2] ),
    .RESET_B(net927),
    .Q(\u_gpio.u_bit[21].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09675_ (.CLK(clknet_1_0__leaf__04479_),
    .D(net34),
    .RESET_B(net921),
    .Q(\u_gpio.u_bit[22].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09676_ (.CLK(clknet_1_0__leaf__04479_),
    .D(net2282),
    .RESET_B(net921),
    .Q(\u_gpio.u_bit[22].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09677_ (.CLK(clknet_1_1__leaf__04479_),
    .D(\u_gpio.u_bit[22].u_dglitch.gpio_ss[1] ),
    .RESET_B(net977),
    .Q(\u_gpio.u_bit[22].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09678_ (.CLK(clknet_1_1__leaf__04479_),
    .D(\u_gpio.u_bit[22].u_dglitch.gpio_ss[2] ),
    .RESET_B(net977),
    .Q(\u_gpio.u_bit[22].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09679_ (.CLK(clknet_1_0__leaf__04480_),
    .D(net1388),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[24].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09680_ (.CLK(clknet_1_1__leaf__04480_),
    .D(net2256),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[24].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09681_ (.CLK(clknet_1_0__leaf__04480_),
    .D(\u_gpio.u_bit[24].u_dglitch.gpio_ss[1] ),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[24].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09682_ (.CLK(clknet_1_1__leaf__04480_),
    .D(\u_gpio.u_bit[24].u_dglitch.gpio_ss[2] ),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[24].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09683_ (.CLK(clknet_1_1__leaf__04481_),
    .D(net36),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[25].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09684_ (.CLK(clknet_1_0__leaf__04481_),
    .D(net2243),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[25].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09685_ (.CLK(clknet_1_1__leaf__04481_),
    .D(\u_gpio.u_bit[25].u_dglitch.gpio_ss[1] ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[25].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09686_ (.CLK(clknet_1_0__leaf__04481_),
    .D(\u_gpio.u_bit[25].u_dglitch.gpio_ss[2] ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[25].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09687_ (.CLK(clknet_1_1__leaf__04482_),
    .D(net1387),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[26].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09688_ (.CLK(clknet_1_0__leaf__04482_),
    .D(net2271),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[26].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09689_ (.CLK(clknet_1_0__leaf__04482_),
    .D(\u_gpio.u_bit[26].u_dglitch.gpio_ss[1] ),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[26].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09690_ (.CLK(clknet_1_1__leaf__04482_),
    .D(\u_gpio.u_bit[26].u_dglitch.gpio_ss[2] ),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[26].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09691_ (.CLK(clknet_1_1__leaf__04483_),
    .D(net38),
    .RESET_B(net850),
    .Q(\u_gpio.u_bit[27].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09692_ (.CLK(clknet_1_1__leaf__04483_),
    .D(net2303),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[27].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09693_ (.CLK(clknet_1_0__leaf__04483_),
    .D(\u_gpio.u_bit[27].u_dglitch.gpio_ss[1] ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[27].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09694_ (.CLK(clknet_1_0__leaf__04483_),
    .D(\u_gpio.u_bit[27].u_dglitch.gpio_ss[2] ),
    .RESET_B(net849),
    .Q(\u_gpio.u_bit[27].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09695_ (.CLK(clknet_1_1__leaf__04484_),
    .D(net4),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[28].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09696_ (.CLK(clknet_1_1__leaf__04484_),
    .D(net2299),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[28].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09697_ (.CLK(clknet_1_0__leaf__04484_),
    .D(\u_gpio.u_bit[28].u_dglitch.gpio_ss[1] ),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[28].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09698_ (.CLK(clknet_1_0__leaf__04484_),
    .D(\u_gpio.u_bit[28].u_dglitch.gpio_ss[2] ),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[28].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09699_ (.CLK(clknet_1_0__leaf__04485_),
    .D(net1306),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[29].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09700_ (.CLK(clknet_1_0__leaf__04485_),
    .D(net2286),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[29].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09701_ (.CLK(clknet_1_1__leaf__04485_),
    .D(\u_gpio.u_bit[29].u_dglitch.gpio_ss[1] ),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[29].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09702_ (.CLK(clknet_1_1__leaf__04485_),
    .D(\u_gpio.u_bit[29].u_dglitch.gpio_ss[2] ),
    .RESET_B(net766),
    .Q(\u_gpio.u_bit[29].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09703_ (.CLK(clknet_1_0__leaf__04486_),
    .D(net24),
    .RESET_B(net875),
    .Q(\u_gpio.u_bit[2].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09704_ (.CLK(clknet_1_1__leaf__04486_),
    .D(net2255),
    .RESET_B(net875),
    .Q(\u_gpio.u_bit[2].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09705_ (.CLK(clknet_1_1__leaf__04486_),
    .D(\u_gpio.u_bit[2].u_dglitch.gpio_ss[1] ),
    .RESET_B(net875),
    .Q(\u_gpio.u_bit[2].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09706_ (.CLK(clknet_1_0__leaf__04486_),
    .D(\u_gpio.u_bit[2].u_dglitch.gpio_ss[2] ),
    .RESET_B(net875),
    .Q(\u_gpio.u_bit[2].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09707_ (.CLK(clknet_1_0__leaf__04487_),
    .D(net1305),
    .RESET_B(net764),
    .Q(\u_gpio.u_bit[30].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09708_ (.CLK(clknet_1_0__leaf__04487_),
    .D(net2300),
    .RESET_B(net764),
    .Q(\u_gpio.u_bit[30].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09709_ (.CLK(clknet_1_1__leaf__04487_),
    .D(\u_gpio.u_bit[30].u_dglitch.gpio_ss[1] ),
    .RESET_B(net764),
    .Q(\u_gpio.u_bit[30].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09710_ (.CLK(clknet_1_1__leaf__04487_),
    .D(\u_gpio.u_bit[30].u_dglitch.gpio_ss[2] ),
    .RESET_B(net763),
    .Q(\u_gpio.u_bit[30].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09711_ (.CLK(clknet_1_0__leaf__04488_),
    .D(net1304),
    .RESET_B(net759),
    .Q(\u_gpio.u_bit[31].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09712_ (.CLK(clknet_1_1__leaf__04488_),
    .D(net2237),
    .RESET_B(net762),
    .Q(\u_gpio.u_bit[31].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09713_ (.CLK(clknet_1_1__leaf__04488_),
    .D(\u_gpio.u_bit[31].u_dglitch.gpio_ss[1] ),
    .RESET_B(net762),
    .Q(\u_gpio.u_bit[31].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09714_ (.CLK(clknet_1_0__leaf__04488_),
    .D(\u_gpio.u_bit[31].u_dglitch.gpio_ss[2] ),
    .RESET_B(net762),
    .Q(\u_gpio.u_bit[31].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09715_ (.CLK(clknet_1_1__leaf__04489_),
    .D(net32),
    .RESET_B(net809),
    .Q(\u_gpio.u_bit[3].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09716_ (.CLK(clknet_1_0__leaf__04489_),
    .D(net2238),
    .RESET_B(net799),
    .Q(\u_gpio.u_bit[3].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09717_ (.CLK(clknet_1_0__leaf__04489_),
    .D(\u_gpio.u_bit[3].u_dglitch.gpio_ss[1] ),
    .RESET_B(net799),
    .Q(\u_gpio.u_bit[3].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09718_ (.CLK(clknet_1_1__leaf__04489_),
    .D(\u_gpio.u_bit[3].u_dglitch.gpio_ss[2] ),
    .RESET_B(net799),
    .Q(\u_gpio.u_bit[3].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09719_ (.CLK(clknet_1_0__leaf__04490_),
    .D(net33),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[4].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09720_ (.CLK(clknet_1_1__leaf__04490_),
    .D(net2249),
    .RESET_B(net880),
    .Q(\u_gpio.u_bit[4].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09721_ (.CLK(clknet_1_0__leaf__04490_),
    .D(\u_gpio.u_bit[4].u_dglitch.gpio_ss[1] ),
    .RESET_B(net881),
    .Q(\u_gpio.u_bit[4].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09722_ (.CLK(clknet_1_1__leaf__04490_),
    .D(\u_gpio.u_bit[4].u_dglitch.gpio_ss[2] ),
    .RESET_B(net881),
    .Q(\u_gpio.u_bit[4].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09723_ (.CLK(clknet_1_0__leaf__04491_),
    .D(net1650),
    .RESET_B(net811),
    .Q(\u_gpio.u_bit[8].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09724_ (.CLK(clknet_1_0__leaf__04491_),
    .D(net2315),
    .RESET_B(net811),
    .Q(\u_gpio.u_bit[8].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09725_ (.CLK(clknet_1_1__leaf__04491_),
    .D(\u_gpio.u_bit[8].u_dglitch.gpio_ss[1] ),
    .RESET_B(net811),
    .Q(\u_gpio.u_bit[8].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09726_ (.CLK(clknet_1_1__leaf__04491_),
    .D(\u_gpio.u_bit[8].u_dglitch.gpio_ss[2] ),
    .RESET_B(net811),
    .Q(\u_gpio.u_bit[8].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09727_ (.CLK(clknet_1_1__leaf__04492_),
    .D(net1571),
    .RESET_B(net798),
    .Q(\u_gpio.u_bit[9].u_dglitch.gpio_ss[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09728_ (.CLK(clknet_1_0__leaf__04492_),
    .D(net2277),
    .RESET_B(net798),
    .Q(\u_gpio.u_bit[9].u_dglitch.gpio_ss[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09729_ (.CLK(clknet_1_0__leaf__04492_),
    .D(\u_gpio.u_bit[9].u_dglitch.gpio_ss[1] ),
    .RESET_B(net800),
    .Q(\u_gpio.u_bit[9].u_dglitch.gpio_ss[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09730_ (.CLK(clknet_1_1__leaf__04492_),
    .D(\u_gpio.u_bit[9].u_dglitch.gpio_ss[2] ),
    .RESET_B(net798),
    .Q(\u_gpio.u_bit[9].u_dglitch.gpio_ss[3] ));
 sky130_fd_sc_hd__dfrtp_4 _09731_ (.CLK(clknet_leaf_21_mclk),
    .D(_00251_),
    .RESET_B(net925),
    .Q(\u_gpio.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _09732_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1815),
    .RESET_B(net976),
    .Q(\u_gpio.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09733_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1846),
    .RESET_B(net977),
    .Q(\u_gpio.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09734_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1819),
    .RESET_B(net979),
    .Q(\u_gpio.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09735_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1833),
    .RESET_B(net977),
    .Q(\u_gpio.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09736_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1821),
    .RESET_B(net977),
    .Q(\u_gpio.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09737_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1830),
    .RESET_B(net978),
    .Q(\u_gpio.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09738_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1849),
    .RESET_B(net811),
    .Q(\u_gpio.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09739_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1838),
    .RESET_B(net799),
    .Q(\u_gpio.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09740_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1869),
    .RESET_B(net814),
    .Q(\u_gpio.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09741_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1852),
    .RESET_B(net923),
    .Q(\u_gpio.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09742_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net2000),
    .RESET_B(net922),
    .Q(\u_gpio.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09743_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1879),
    .RESET_B(net802),
    .Q(\u_gpio.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09744_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1900),
    .RESET_B(net802),
    .Q(\u_gpio.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09745_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1896),
    .RESET_B(net802),
    .Q(\u_gpio.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09746_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1936),
    .RESET_B(net915),
    .Q(\u_gpio.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09747_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1954),
    .RESET_B(net916),
    .Q(\u_gpio.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09748_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1862),
    .RESET_B(net923),
    .Q(\u_gpio.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09749_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1958),
    .RESET_B(net923),
    .Q(\u_gpio.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09750_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1952),
    .RESET_B(net920),
    .Q(\u_gpio.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09751_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1947),
    .RESET_B(net926),
    .Q(\u_gpio.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09752_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1942),
    .RESET_B(net919),
    .Q(\u_gpio.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09753_ (.CLK(clknet_2_2__leaf__04493_),
    .D(net1956),
    .RESET_B(net925),
    .Q(\u_gpio.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09754_ (.CLK(clknet_2_3__leaf__04493_),
    .D(net1963),
    .RESET_B(net923),
    .Q(\u_gpio.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09755_ (.CLK(clknet_2_2__leaf__04493_),
    .D(\u_gpio.u_reg.reg_out[23] ),
    .RESET_B(net918),
    .Q(\u_gpio.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09756_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1950),
    .RESET_B(net799),
    .Q(\u_gpio.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09757_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1925),
    .RESET_B(net796),
    .Q(\u_gpio.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09758_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1938),
    .RESET_B(net796),
    .Q(\u_gpio.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09759_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1911),
    .RESET_B(net852),
    .Q(\u_gpio.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09760_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1842),
    .RESET_B(net796),
    .Q(\u_gpio.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09761_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1945),
    .RESET_B(net798),
    .Q(\u_gpio.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09762_ (.CLK(clknet_2_0__leaf__04493_),
    .D(net1981),
    .RESET_B(net798),
    .Q(\u_gpio.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09763_ (.CLK(clknet_2_1__leaf__04493_),
    .D(net1921),
    .RESET_B(net796),
    .Q(\u_gpio.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09764_ (.CLK(clknet_1_0__leaf__04546_),
    .D(net1607),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09765_ (.CLK(clknet_1_1__leaf__04546_),
    .D(net1600),
    .RESET_B(net925),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09766_ (.CLK(clknet_1_0__leaf__04546_),
    .D(net1589),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09767_ (.CLK(clknet_1_1__leaf__04546_),
    .D(net1582),
    .RESET_B(net927),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09768_ (.CLK(clknet_1_0__leaf__04546_),
    .D(net1567),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09769_ (.CLK(clknet_1_1__leaf__04546_),
    .D(net1559),
    .RESET_B(net927),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09770_ (.CLK(clknet_1_0__leaf__04546_),
    .D(net1552),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09771_ (.CLK(clknet_1_1__leaf__04546_),
    .D(net1545),
    .RESET_B(net919),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09772_ (.CLK(clknet_1_0__leaf__04547_),
    .D(net1536),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09773_ (.CLK(clknet_1_1__leaf__04547_),
    .D(net1528),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09774_ (.CLK(clknet_1_1__leaf__04547_),
    .D(net1521),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09775_ (.CLK(clknet_1_1__leaf__04547_),
    .D(net1514),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09776_ (.CLK(clknet_1_1__leaf__04547_),
    .D(net1507),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09777_ (.CLK(clknet_1_0__leaf__04547_),
    .D(net1499),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09778_ (.CLK(clknet_1_0__leaf__04547_),
    .D(net1483),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09779_ (.CLK(clknet_1_0__leaf__04547_),
    .D(net1476),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09780_ (.CLK(clknet_1_1__leaf__04548_),
    .D(net1296),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09781_ (.CLK(clknet_1_0__leaf__04548_),
    .D(net1575),
    .RESET_B(net857),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09782_ (.CLK(clknet_1_1__leaf__04548_),
    .D(net1490),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09783_ (.CLK(clknet_1_0__leaf__04548_),
    .D(net1467),
    .RESET_B(net868),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09784_ (.CLK(clknet_1_0__leaf__04548_),
    .D(net1460),
    .RESET_B(net856),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09785_ (.CLK(clknet_1_1__leaf__04548_),
    .D(net1450),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09786_ (.CLK(clknet_1_1__leaf__04548_),
    .D(net1444),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09787_ (.CLK(clknet_1_0__leaf__04548_),
    .D(net1436),
    .RESET_B(net858),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09788_ (.CLK(clknet_1_1__leaf__04549_),
    .D(net1426),
    .RESET_B(net811),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09789_ (.CLK(clknet_1_0__leaf__04549_),
    .D(net1420),
    .RESET_B(net800),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09790_ (.CLK(clknet_1_0__leaf__04549_),
    .D(net1287),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09791_ (.CLK(clknet_1_0__leaf__04549_),
    .D(net1643),
    .RESET_B(net792),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09792_ (.CLK(clknet_1_0__leaf__04549_),
    .D(net1637),
    .RESET_B(net808),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09793_ (.CLK(clknet_1_1__leaf__04549_),
    .D(net1629),
    .RESET_B(net804),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09794_ (.CLK(clknet_1_1__leaf__04549_),
    .D(net1622),
    .RESET_B(net804),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09795_ (.CLK(clknet_1_1__leaf__04549_),
    .D(net1614),
    .RESET_B(net806),
    .Q(\u_gpio.cfg_gpio_negedge_int_sel[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09796_ (.CLK(clknet_1_0__leaf__04542_),
    .D(net1607),
    .RESET_B(net923),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09797_ (.CLK(clknet_1_1__leaf__04542_),
    .D(net1600),
    .RESET_B(net930),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09798_ (.CLK(clknet_1_0__leaf__04542_),
    .D(net1589),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09799_ (.CLK(clknet_1_1__leaf__04542_),
    .D(net1581),
    .RESET_B(net926),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09800_ (.CLK(clknet_1_1__leaf__04542_),
    .D(net1567),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09801_ (.CLK(clknet_1_1__leaf__04542_),
    .D(net1559),
    .RESET_B(net926),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09802_ (.CLK(clknet_1_0__leaf__04542_),
    .D(net1552),
    .RESET_B(net923),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09803_ (.CLK(clknet_1_0__leaf__04542_),
    .D(net1545),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09804_ (.CLK(clknet_1_0__leaf__04543_),
    .D(net1536),
    .RESET_B(net766),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09805_ (.CLK(clknet_1_1__leaf__04543_),
    .D(net1528),
    .RESET_B(net767),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09806_ (.CLK(clknet_1_1__leaf__04543_),
    .D(net1521),
    .RESET_B(net767),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09807_ (.CLK(clknet_1_1__leaf__04543_),
    .D(net1514),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09808_ (.CLK(clknet_1_1__leaf__04543_),
    .D(net1507),
    .RESET_B(net769),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09809_ (.CLK(clknet_1_0__leaf__04543_),
    .D(net1499),
    .RESET_B(net768),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09810_ (.CLK(clknet_1_0__leaf__04543_),
    .D(net1483),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09811_ (.CLK(clknet_1_0__leaf__04543_),
    .D(net1476),
    .RESET_B(net770),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09812_ (.CLK(clknet_1_1__leaf__04544_),
    .D(net1296),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09813_ (.CLK(clknet_1_0__leaf__04544_),
    .D(net1575),
    .RESET_B(net857),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09814_ (.CLK(clknet_1_1__leaf__04544_),
    .D(net1490),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09815_ (.CLK(clknet_1_0__leaf__04544_),
    .D(net1467),
    .RESET_B(net868),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09816_ (.CLK(clknet_1_0__leaf__04544_),
    .D(net1460),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09817_ (.CLK(clknet_1_1__leaf__04544_),
    .D(net1450),
    .RESET_B(net871),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09818_ (.CLK(clknet_1_1__leaf__04544_),
    .D(net1444),
    .RESET_B(net869),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09819_ (.CLK(clknet_1_0__leaf__04544_),
    .D(net1436),
    .RESET_B(net858),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09820_ (.CLK(clknet_1_1__leaf__04545_),
    .D(net1426),
    .RESET_B(net811),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09821_ (.CLK(clknet_1_0__leaf__04545_),
    .D(net1420),
    .RESET_B(net808),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09822_ (.CLK(clknet_1_0__leaf__04545_),
    .D(net1287),
    .RESET_B(net802),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09823_ (.CLK(clknet_1_0__leaf__04545_),
    .D(net1643),
    .RESET_B(net801),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09824_ (.CLK(clknet_1_0__leaf__04545_),
    .D(net1637),
    .RESET_B(net803),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09825_ (.CLK(clknet_1_1__leaf__04545_),
    .D(net1629),
    .RESET_B(net801),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09826_ (.CLK(clknet_1_1__leaf__04545_),
    .D(net1622),
    .RESET_B(net804),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09827_ (.CLK(clknet_1_1__leaf__04545_),
    .D(net1614),
    .RESET_B(net806),
    .Q(\u_gpio.cfg_gpio_posedge_int_sel[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09828_ (.CLK(clknet_1_0__leaf__04538_),
    .D(net1606),
    .RESET_B(net919),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09829_ (.CLK(clknet_1_1__leaf__04538_),
    .D(net1599),
    .RESET_B(net925),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09830_ (.CLK(clknet_1_0__leaf__04538_),
    .D(net1590),
    .RESET_B(net917),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09831_ (.CLK(clknet_1_1__leaf__04538_),
    .D(net1581),
    .RESET_B(net926),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09832_ (.CLK(clknet_1_1__leaf__04538_),
    .D(net1567),
    .RESET_B(net917),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09833_ (.CLK(clknet_1_1__leaf__04538_),
    .D(net1560),
    .RESET_B(net926),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09834_ (.CLK(clknet_1_0__leaf__04538_),
    .D(net1550),
    .RESET_B(net918),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09835_ (.CLK(clknet_1_0__leaf__04538_),
    .D(net1545),
    .RESET_B(net918),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09836_ (.CLK(clknet_1_0__leaf__04539_),
    .D(net1537),
    .RESET_B(net795),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09837_ (.CLK(clknet_1_1__leaf__04539_),
    .D(net1529),
    .RESET_B(net771),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09838_ (.CLK(clknet_1_1__leaf__04539_),
    .D(net1522),
    .RESET_B(net771),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09839_ (.CLK(clknet_1_1__leaf__04539_),
    .D(net1514),
    .RESET_B(net769),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09840_ (.CLK(clknet_1_1__leaf__04539_),
    .D(net1507),
    .RESET_B(net796),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09841_ (.CLK(clknet_1_0__leaf__04539_),
    .D(net1499),
    .RESET_B(net795),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09842_ (.CLK(clknet_1_0__leaf__04539_),
    .D(net1485),
    .RESET_B(net770),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09843_ (.CLK(clknet_1_0__leaf__04539_),
    .D(net1477),
    .RESET_B(net770),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09844_ (.CLK(clknet_1_1__leaf__04540_),
    .D(net1296),
    .RESET_B(net869),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09845_ (.CLK(clknet_1_0__leaf__04540_),
    .D(net1574),
    .RESET_B(net857),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09846_ (.CLK(clknet_1_1__leaf__04540_),
    .D(net1490),
    .RESET_B(net869),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09847_ (.CLK(clknet_1_0__leaf__04540_),
    .D(net1468),
    .RESET_B(net868),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09848_ (.CLK(clknet_1_0__leaf__04540_),
    .D(net1460),
    .RESET_B(net868),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09849_ (.CLK(clknet_1_1__leaf__04540_),
    .D(net1450),
    .RESET_B(net869),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09850_ (.CLK(clknet_1_1__leaf__04540_),
    .D(net1444),
    .RESET_B(net869),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09851_ (.CLK(clknet_1_0__leaf__04540_),
    .D(net1436),
    .RESET_B(net857),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09852_ (.CLK(clknet_1_1__leaf__04541_),
    .D(net1426),
    .RESET_B(net805),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09853_ (.CLK(clknet_1_0__leaf__04541_),
    .D(net1420),
    .RESET_B(net802),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09854_ (.CLK(clknet_1_0__leaf__04541_),
    .D(net1287),
    .RESET_B(net802),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09855_ (.CLK(clknet_1_0__leaf__04541_),
    .D(net1643),
    .RESET_B(net801),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09856_ (.CLK(clknet_1_0__leaf__04541_),
    .D(net1637),
    .RESET_B(net802),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09857_ (.CLK(clknet_1_1__leaf__04541_),
    .D(net1629),
    .RESET_B(net804),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09858_ (.CLK(clknet_1_1__leaf__04541_),
    .D(net1622),
    .RESET_B(net804),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09859_ (.CLK(clknet_1_1__leaf__04541_),
    .D(net1614),
    .RESET_B(net805),
    .Q(\u_gpio.u_reg.cfg_gpio_int_mask[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09860_ (.CLK(_04506_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .RESET_B(net870),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09861_ (.CLK(_04507_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.hware_req ),
    .RESET_B(net793),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[10].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09862_ (.CLK(_04508_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.hware_req ),
    .RESET_B(net792),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09863_ (.CLK(_04509_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.hware_req ),
    .RESET_B(net802),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09864_ (.CLK(_04510_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.hware_req ),
    .RESET_B(net801),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09865_ (.CLK(_04511_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.hware_req ),
    .RESET_B(net804),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[14].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09866_ (.CLK(_04512_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.hware_req ),
    .RESET_B(net916),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09867_ (.CLK(_04513_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.hware_req ),
    .RESET_B(net923),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09868_ (.CLK(_04514_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.hware_req ),
    .RESET_B(net918),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09869_ (.CLK(_04515_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.hware_req ),
    .RESET_B(net915),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09870_ (.CLK(_04516_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.hware_req ),
    .RESET_B(net926),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09871_ (.CLK(_04517_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .RESET_B(net857),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09872_ (.CLK(_04518_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.hware_req ),
    .RESET_B(net917),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09873_ (.CLK(_04519_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.hware_req ),
    .RESET_B(net926),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09874_ (.CLK(_04520_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.hware_req ),
    .RESET_B(net922),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09875_ (.CLK(_04521_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.hware_req ),
    .RESET_B(net915),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09876_ (.CLK(_04522_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.hware_req ),
    .RESET_B(net768),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09877_ (.CLK(_04523_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.hware_req ),
    .RESET_B(net767),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[25].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09878_ (.CLK(_04524_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.hware_req ),
    .RESET_B(net767),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09879_ (.CLK(_04525_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.hware_req ),
    .RESET_B(net769),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09880_ (.CLK(_04526_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.hware_req ),
    .RESET_B(net796),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09881_ (.CLK(_04527_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.hware_req ),
    .RESET_B(net768),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09882_ (.CLK(_04528_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .RESET_B(net870),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09883_ (.CLK(_04529_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.hware_req ),
    .RESET_B(net764),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[30].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09884_ (.CLK(_04530_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.hware_req ),
    .RESET_B(net770),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09885_ (.CLK(_04531_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.hware_req ),
    .RESET_B(net868),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[3].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09886_ (.CLK(_04532_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.hware_req ),
    .RESET_B(net867),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09887_ (.CLK(_04533_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.hware_req ),
    .RESET_B(net869),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09888_ (.CLK(_04534_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.hware_req ),
    .RESET_B(net868),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09889_ (.CLK(_04535_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.hware_req ),
    .RESET_B(net856),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09890_ (.CLK(_04536_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.hware_req ),
    .RESET_B(net811),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09891_ (.CLK(_04537_),
    .D(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.hware_req ),
    .RESET_B(net808),
    .Q(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _09892_ (.CLK(clknet_1_1__leaf__04502_),
    .D(net1607),
    .RESET_B(net925),
    .Q(\u_gpio.cfg_gpio_out_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09893_ (.CLK(clknet_1_1__leaf__04502_),
    .D(net1600),
    .RESET_B(net925),
    .Q(\u_gpio.cfg_gpio_out_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09894_ (.CLK(clknet_1_0__leaf__04502_),
    .D(net1590),
    .RESET_B(net904),
    .Q(\u_gpio.cfg_gpio_out_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09895_ (.CLK(clknet_1_0__leaf__04502_),
    .D(net1581),
    .RESET_B(net910),
    .Q(\u_gpio.cfg_gpio_out_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09896_ (.CLK(clknet_1_0__leaf__04502_),
    .D(net1567),
    .RESET_B(net910),
    .Q(\u_gpio.cfg_gpio_out_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09897_ (.CLK(clknet_1_0__leaf__04502_),
    .D(net1560),
    .RESET_B(net910),
    .Q(\u_gpio.cfg_gpio_out_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09898_ (.CLK(clknet_1_1__leaf__04502_),
    .D(net1552),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_out_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09899_ (.CLK(clknet_1_1__leaf__04502_),
    .D(net1545),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_out_data[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09900_ (.CLK(clknet_1_0__leaf__04503_),
    .D(net1537),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_data[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09901_ (.CLK(clknet_1_1__leaf__04503_),
    .D(net1529),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_data[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09902_ (.CLK(clknet_1_1__leaf__04503_),
    .D(net1522),
    .RESET_B(net796),
    .Q(\u_gpio.cfg_gpio_out_data[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09903_ (.CLK(clknet_1_1__leaf__04503_),
    .D(net1516),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_out_data[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09904_ (.CLK(clknet_1_1__leaf__04503_),
    .D(net1508),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_out_data[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09905_ (.CLK(clknet_1_0__leaf__04503_),
    .D(net1500),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_out_data[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09906_ (.CLK(clknet_1_0__leaf__04503_),
    .D(net1484),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_data[30] ));
 sky130_fd_sc_hd__dfrtp_1 _09907_ (.CLK(clknet_1_0__leaf__04503_),
    .D(net1478),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_data[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09908_ (.CLK(clknet_1_1__leaf__04504_),
    .D(net1296),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_out_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09909_ (.CLK(clknet_1_0__leaf__04504_),
    .D(net1574),
    .RESET_B(net857),
    .Q(\u_gpio.cfg_gpio_out_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09910_ (.CLK(clknet_1_1__leaf__04504_),
    .D(net1490),
    .RESET_B(net869),
    .Q(\u_gpio.cfg_gpio_out_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09911_ (.CLK(clknet_1_0__leaf__04504_),
    .D(net1468),
    .RESET_B(net868),
    .Q(\u_gpio.cfg_gpio_out_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09912_ (.CLK(clknet_1_0__leaf__04504_),
    .D(net1460),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_out_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09913_ (.CLK(clknet_1_1__leaf__04504_),
    .D(net1450),
    .RESET_B(net869),
    .Q(\u_gpio.cfg_gpio_out_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09914_ (.CLK(clknet_1_1__leaf__04504_),
    .D(net1444),
    .RESET_B(net869),
    .Q(\u_gpio.cfg_gpio_out_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09915_ (.CLK(clknet_1_0__leaf__04504_),
    .D(net1436),
    .RESET_B(net856),
    .Q(\u_gpio.cfg_gpio_out_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09916_ (.CLK(clknet_1_1__leaf__04505_),
    .D(net1426),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_out_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09917_ (.CLK(clknet_1_0__leaf__04505_),
    .D(net1420),
    .RESET_B(net802),
    .Q(\u_gpio.cfg_gpio_out_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09918_ (.CLK(clknet_1_0__leaf__04505_),
    .D(net1287),
    .RESET_B(net794),
    .Q(\u_gpio.cfg_gpio_out_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09919_ (.CLK(clknet_1_0__leaf__04505_),
    .D(net1643),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_out_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09920_ (.CLK(clknet_1_0__leaf__04505_),
    .D(net1637),
    .RESET_B(net802),
    .Q(\u_gpio.cfg_gpio_out_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09921_ (.CLK(clknet_1_1__leaf__04505_),
    .D(net1629),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_out_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09922_ (.CLK(clknet_1_1__leaf__04505_),
    .D(net1622),
    .RESET_B(net806),
    .Q(\u_gpio.cfg_gpio_out_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09923_ (.CLK(clknet_1_1__leaf__04505_),
    .D(net1615),
    .RESET_B(net806),
    .Q(\u_gpio.cfg_gpio_out_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09924_ (.CLK(clknet_1_0__leaf__04498_),
    .D(net1606),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_out_type[16] ));
 sky130_fd_sc_hd__dfrtp_1 _09925_ (.CLK(clknet_1_1__leaf__04498_),
    .D(net1599),
    .RESET_B(net925),
    .Q(\u_gpio.cfg_gpio_out_type[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09926_ (.CLK(clknet_1_0__leaf__04498_),
    .D(net1590),
    .RESET_B(net905),
    .Q(\u_gpio.cfg_gpio_out_type[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09927_ (.CLK(clknet_1_1__leaf__04498_),
    .D(net1581),
    .RESET_B(net926),
    .Q(\u_gpio.cfg_gpio_out_type[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09928_ (.CLK(clknet_1_1__leaf__04498_),
    .D(net1567),
    .RESET_B(net904),
    .Q(\u_gpio.cfg_gpio_out_type[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09929_ (.CLK(clknet_1_1__leaf__04498_),
    .D(net1560),
    .RESET_B(net926),
    .Q(\u_gpio.cfg_gpio_out_type[21] ));
 sky130_fd_sc_hd__dfrtp_2 _09930_ (.CLK(clknet_1_0__leaf__04498_),
    .D(net1552),
    .RESET_B(net918),
    .Q(\u_gpio.cfg_gpio_out_type[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09931_ (.CLK(clknet_1_0__leaf__04498_),
    .D(net1545),
    .RESET_B(net917),
    .Q(\u_gpio.cfg_gpio_out_type[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09932_ (.CLK(clknet_1_0__leaf__04499_),
    .D(net1538),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_type[24] ));
 sky130_fd_sc_hd__dfrtp_2 _09933_ (.CLK(clknet_1_1__leaf__04499_),
    .D(net1530),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_out_type[25] ));
 sky130_fd_sc_hd__dfrtp_2 _09934_ (.CLK(clknet_1_1__leaf__04499_),
    .D(net1523),
    .RESET_B(net796),
    .Q(\u_gpio.cfg_gpio_out_type[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09935_ (.CLK(clknet_1_1__leaf__04499_),
    .D(net1516),
    .RESET_B(net799),
    .Q(\u_gpio.cfg_gpio_out_type[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09936_ (.CLK(clknet_1_1__leaf__04499_),
    .D(net1508),
    .RESET_B(net799),
    .Q(\u_gpio.cfg_gpio_out_type[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09937_ (.CLK(clknet_1_0__leaf__04499_),
    .D(net1500),
    .RESET_B(net798),
    .Q(\u_gpio.cfg_gpio_out_type[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09938_ (.CLK(clknet_1_0__leaf__04499_),
    .D(net1484),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_out_type[30] ));
 sky130_fd_sc_hd__dfrtp_4 _09939_ (.CLK(clknet_1_0__leaf__04499_),
    .D(net1478),
    .RESET_B(net798),
    .Q(\u_gpio.cfg_gpio_out_type[31] ));
 sky130_fd_sc_hd__dfrtp_1 _09940_ (.CLK(clknet_1_1__leaf__04500_),
    .D(net1296),
    .RESET_B(net870),
    .Q(\u_gpio.cfg_gpio_out_type[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09941_ (.CLK(clknet_1_0__leaf__04500_),
    .D(net1574),
    .RESET_B(net857),
    .Q(\u_gpio.cfg_gpio_out_type[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09942_ (.CLK(clknet_1_1__leaf__04500_),
    .D(net1490),
    .RESET_B(net871),
    .Q(\u_gpio.cfg_gpio_out_type[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09943_ (.CLK(clknet_1_0__leaf__04500_),
    .D(net1468),
    .RESET_B(net868),
    .Q(\u_gpio.cfg_gpio_out_type[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09944_ (.CLK(clknet_1_0__leaf__04500_),
    .D(net1460),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_out_type[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09945_ (.CLK(clknet_1_1__leaf__04500_),
    .D(net1450),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_out_type[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09946_ (.CLK(clknet_1_1__leaf__04500_),
    .D(net1444),
    .RESET_B(net869),
    .Q(\u_gpio.cfg_gpio_out_type[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09947_ (.CLK(clknet_1_0__leaf__04500_),
    .D(net1436),
    .RESET_B(net856),
    .Q(\u_gpio.cfg_gpio_out_type[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09948_ (.CLK(clknet_1_1__leaf__04501_),
    .D(net1426),
    .RESET_B(net922),
    .Q(\u_gpio.cfg_gpio_out_type[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09949_ (.CLK(clknet_1_0__leaf__04501_),
    .D(net1420),
    .RESET_B(net808),
    .Q(\u_gpio.cfg_gpio_out_type[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09950_ (.CLK(clknet_1_0__leaf__04501_),
    .D(net1287),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_out_type[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09951_ (.CLK(clknet_1_0__leaf__04501_),
    .D(net1643),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_out_type[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09952_ (.CLK(clknet_1_1__leaf__04501_),
    .D(net1637),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_out_type[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09953_ (.CLK(clknet_1_0__leaf__04501_),
    .D(net1629),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_out_type[13] ));
 sky130_fd_sc_hd__dfrtp_2 _09954_ (.CLK(clknet_1_1__leaf__04501_),
    .D(net1622),
    .RESET_B(net806),
    .Q(\u_gpio.cfg_gpio_out_type[14] ));
 sky130_fd_sc_hd__dfrtp_2 _09955_ (.CLK(clknet_1_1__leaf__04501_),
    .D(net1615),
    .RESET_B(net915),
    .Q(\u_gpio.cfg_gpio_out_type[15] ));
 sky130_fd_sc_hd__dfrtp_4 _09956_ (.CLK(clknet_1_1__leaf__04494_),
    .D(net1607),
    .RESET_B(net925),
    .Q(\u_gpio.cfg_gpio_dir_sel[16] ));
 sky130_fd_sc_hd__dfrtp_4 _09957_ (.CLK(clknet_1_1__leaf__04494_),
    .D(net1599),
    .RESET_B(net929),
    .Q(\u_gpio.cfg_gpio_dir_sel[17] ));
 sky130_fd_sc_hd__dfrtp_1 _09958_ (.CLK(clknet_1_0__leaf__04494_),
    .D(net1590),
    .RESET_B(net905),
    .Q(\u_gpio.cfg_gpio_dir_sel[18] ));
 sky130_fd_sc_hd__dfrtp_1 _09959_ (.CLK(clknet_1_0__leaf__04494_),
    .D(net1581),
    .RESET_B(net911),
    .Q(\u_gpio.cfg_gpio_dir_sel[19] ));
 sky130_fd_sc_hd__dfrtp_1 _09960_ (.CLK(clknet_1_0__leaf__04494_),
    .D(net1567),
    .RESET_B(net910),
    .Q(\u_gpio.cfg_gpio_dir_sel[20] ));
 sky130_fd_sc_hd__dfrtp_1 _09961_ (.CLK(clknet_1_0__leaf__04494_),
    .D(net1560),
    .RESET_B(net911),
    .Q(\u_gpio.cfg_gpio_dir_sel[21] ));
 sky130_fd_sc_hd__dfrtp_1 _09962_ (.CLK(clknet_1_1__leaf__04494_),
    .D(net1553),
    .RESET_B(net919),
    .Q(\u_gpio.cfg_gpio_dir_sel[22] ));
 sky130_fd_sc_hd__dfrtp_1 _09963_ (.CLK(clknet_1_1__leaf__04494_),
    .D(net1547),
    .RESET_B(net919),
    .Q(\u_gpio.cfg_gpio_dir_sel[23] ));
 sky130_fd_sc_hd__dfrtp_1 _09964_ (.CLK(clknet_1_1__leaf__04495_),
    .D(net1538),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_dir_sel[24] ));
 sky130_fd_sc_hd__dfrtp_1 _09965_ (.CLK(clknet_1_0__leaf__04495_),
    .D(net1530),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_dir_sel[25] ));
 sky130_fd_sc_hd__dfrtp_1 _09966_ (.CLK(clknet_1_0__leaf__04495_),
    .D(net1523),
    .RESET_B(net797),
    .Q(\u_gpio.cfg_gpio_dir_sel[26] ));
 sky130_fd_sc_hd__dfrtp_1 _09967_ (.CLK(clknet_1_0__leaf__04495_),
    .D(net1516),
    .RESET_B(net796),
    .Q(\u_gpio.cfg_gpio_dir_sel[27] ));
 sky130_fd_sc_hd__dfrtp_1 _09968_ (.CLK(clknet_1_1__leaf__04495_),
    .D(net1508),
    .RESET_B(net799),
    .Q(\u_gpio.cfg_gpio_dir_sel[28] ));
 sky130_fd_sc_hd__dfrtp_1 _09969_ (.CLK(clknet_1_1__leaf__04495_),
    .D(net1500),
    .RESET_B(net798),
    .Q(\u_gpio.cfg_gpio_dir_sel[29] ));
 sky130_fd_sc_hd__dfrtp_1 _09970_ (.CLK(clknet_1_0__leaf__04495_),
    .D(net1484),
    .RESET_B(net795),
    .Q(\u_gpio.cfg_gpio_dir_sel[30] ));
 sky130_fd_sc_hd__dfrtp_4 _09971_ (.CLK(clknet_1_1__leaf__04495_),
    .D(net1478),
    .RESET_B(net798),
    .Q(\u_gpio.cfg_gpio_dir_sel[31] ));
 sky130_fd_sc_hd__dfrtp_2 _09972_ (.CLK(clknet_1_1__leaf__04496_),
    .D(net1296),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_dir_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09973_ (.CLK(clknet_1_0__leaf__04496_),
    .D(net1574),
    .RESET_B(net856),
    .Q(\u_gpio.cfg_gpio_dir_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09974_ (.CLK(clknet_1_0__leaf__04496_),
    .D(net1490),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_dir_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09975_ (.CLK(clknet_1_0__leaf__04496_),
    .D(net1468),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_dir_sel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09976_ (.CLK(clknet_1_1__leaf__04496_),
    .D(net1461),
    .RESET_B(net867),
    .Q(\u_gpio.cfg_gpio_dir_sel[4] ));
 sky130_fd_sc_hd__dfrtp_1 _09977_ (.CLK(clknet_1_1__leaf__04496_),
    .D(net1450),
    .RESET_B(net871),
    .Q(\u_gpio.cfg_gpio_dir_sel[5] ));
 sky130_fd_sc_hd__dfrtp_1 _09978_ (.CLK(clknet_1_1__leaf__04496_),
    .D(net1444),
    .RESET_B(net868),
    .Q(\u_gpio.cfg_gpio_dir_sel[6] ));
 sky130_fd_sc_hd__dfrtp_1 _09979_ (.CLK(clknet_1_0__leaf__04496_),
    .D(net1436),
    .RESET_B(net858),
    .Q(\u_gpio.cfg_gpio_dir_sel[7] ));
 sky130_fd_sc_hd__dfrtp_1 _09980_ (.CLK(clknet_1_1__leaf__04497_),
    .D(net1426),
    .RESET_B(net922),
    .Q(\u_gpio.cfg_gpio_dir_sel[8] ));
 sky130_fd_sc_hd__dfrtp_1 _09981_ (.CLK(clknet_1_0__leaf__04497_),
    .D(net1422),
    .RESET_B(net800),
    .Q(\u_gpio.cfg_gpio_dir_sel[9] ));
 sky130_fd_sc_hd__dfrtp_1 _09982_ (.CLK(clknet_1_0__leaf__04497_),
    .D(net1287),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_dir_sel[10] ));
 sky130_fd_sc_hd__dfrtp_1 _09983_ (.CLK(clknet_1_0__leaf__04497_),
    .D(net1644),
    .RESET_B(net793),
    .Q(\u_gpio.cfg_gpio_dir_sel[11] ));
 sky130_fd_sc_hd__dfrtp_1 _09984_ (.CLK(clknet_1_1__leaf__04497_),
    .D(net1637),
    .RESET_B(net811),
    .Q(\u_gpio.cfg_gpio_dir_sel[12] ));
 sky130_fd_sc_hd__dfrtp_1 _09985_ (.CLK(clknet_1_0__leaf__04497_),
    .D(net1629),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_dir_sel[13] ));
 sky130_fd_sc_hd__dfrtp_1 _09986_ (.CLK(clknet_1_1__leaf__04497_),
    .D(net1622),
    .RESET_B(net805),
    .Q(\u_gpio.cfg_gpio_dir_sel[14] ));
 sky130_fd_sc_hd__dfrtp_1 _09987_ (.CLK(clknet_1_1__leaf__04497_),
    .D(net1615),
    .RESET_B(net916),
    .Q(\u_gpio.cfg_gpio_dir_sel[15] ));
 sky130_fd_sc_hd__dfrtp_1 _09988_ (.CLK(\u_glbl_reg.dbg_clk_ref_buf ),
    .D(_00043_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.dbg_clk_div16 ));
 sky130_fd_sc_hd__dfrtp_1 _09989_ (.CLK(clknet_1_1__leaf__04355_),
    .D(_00046_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.low_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09990_ (.CLK(clknet_1_0__leaf__04355_),
    .D(_00047_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.low_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09991_ (.CLK(clknet_1_0__leaf__04355_),
    .D(_00048_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.low_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09992_ (.CLK(clknet_1_1__leaf__04355_),
    .D(_00049_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.low_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _09993_ (.CLK(clknet_1_0__leaf__04354_),
    .D(_00039_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.high_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09994_ (.CLK(clknet_1_0__leaf__04354_),
    .D(_00040_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.high_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _09995_ (.CLK(clknet_1_1__leaf__04354_),
    .D(_00041_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.high_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _09996_ (.CLK(clknet_1_1__leaf__04354_),
    .D(_00042_),
    .RESET_B(net1386),
    .Q(\u_glbl_reg.u_dbgclk.high_count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _09997_ (.CLK(clknet_1_1__leaf_user_clock1),
    .D(_00053_),
    .RESET_B(net1380),
    .Q(net365));
 sky130_fd_sc_hd__dfrtp_1 _09998_ (.CLK(clknet_1_1__leaf__04357_),
    .D(_00056_),
    .RESET_B(net1380),
    .Q(\u_glbl_reg.u_pll_ref_clk.low_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _09999_ (.CLK(clknet_1_0__leaf__04357_),
    .D(_00057_),
    .RESET_B(net1380),
    .Q(\u_glbl_reg.u_pll_ref_clk.low_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10000_ (.CLK(clknet_1_0__leaf__04357_),
    .D(_00058_),
    .RESET_B(net1380),
    .Q(\u_glbl_reg.u_pll_ref_clk.low_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10001_ (.CLK(clknet_1_0__leaf__04356_),
    .D(_00050_),
    .RESET_B(net1381),
    .Q(\u_glbl_reg.u_pll_ref_clk.high_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10002_ (.CLK(clknet_1_0__leaf__04356_),
    .D(_00051_),
    .RESET_B(net1381),
    .Q(\u_glbl_reg.u_pll_ref_clk.high_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10003_ (.CLK(clknet_1_1__leaf__04356_),
    .D(_00052_),
    .RESET_B(net1381),
    .Q(\u_glbl_reg.u_pll_ref_clk.high_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10004_ (.CLK(clknet_leaf_23_mclk),
    .D(_00702_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10005_ (.CLK(clknet_leaf_23_mclk),
    .D(_00713_),
    .RESET_B(net914),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10006_ (.CLK(clknet_leaf_32_mclk),
    .D(_00724_),
    .RESET_B(net911),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10007_ (.CLK(clknet_leaf_31_mclk),
    .D(_00727_),
    .RESET_B(net912),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10008_ (.CLK(clknet_leaf_32_mclk),
    .D(_00728_),
    .RESET_B(net912),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10009_ (.CLK(clknet_leaf_31_mclk),
    .D(_00729_),
    .RESET_B(net912),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10010_ (.CLK(clknet_leaf_31_mclk),
    .D(_00730_),
    .RESET_B(net912),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10011_ (.CLK(clknet_leaf_31_mclk),
    .D(_00731_),
    .RESET_B(net908),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10012_ (.CLK(clknet_leaf_31_mclk),
    .D(_00732_),
    .RESET_B(net908),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10013_ (.CLK(clknet_leaf_31_mclk),
    .D(_00733_),
    .RESET_B(net914),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10014_ (.CLK(clknet_leaf_31_mclk),
    .D(_00703_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10015_ (.CLK(clknet_leaf_30_mclk),
    .D(_00704_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10016_ (.CLK(clknet_leaf_30_mclk),
    .D(_00705_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10017_ (.CLK(clknet_leaf_30_mclk),
    .D(_00706_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10018_ (.CLK(clknet_leaf_30_mclk),
    .D(_00707_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10019_ (.CLK(clknet_leaf_33_mclk),
    .D(_00708_),
    .RESET_B(net943),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10020_ (.CLK(clknet_leaf_43_mclk),
    .D(_00709_),
    .RESET_B(net943),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10021_ (.CLK(clknet_leaf_43_mclk),
    .D(_00710_),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10022_ (.CLK(clknet_leaf_43_mclk),
    .D(_00711_),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10023_ (.CLK(clknet_leaf_43_mclk),
    .D(_00712_),
    .RESET_B(net945),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10024_ (.CLK(clknet_leaf_33_mclk),
    .D(_00714_),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10025_ (.CLK(clknet_leaf_33_mclk),
    .D(_00715_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10026_ (.CLK(clknet_leaf_32_mclk),
    .D(_00716_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10027_ (.CLK(clknet_leaf_33_mclk),
    .D(_00717_),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10028_ (.CLK(clknet_leaf_32_mclk),
    .D(_00718_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10029_ (.CLK(clknet_leaf_32_mclk),
    .D(_00719_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10030_ (.CLK(clknet_leaf_32_mclk),
    .D(_00720_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10031_ (.CLK(clknet_leaf_31_mclk),
    .D(_00721_),
    .RESET_B(net913),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10032_ (.CLK(clknet_leaf_31_mclk),
    .D(_00722_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10033_ (.CLK(clknet_leaf_31_mclk),
    .D(_00723_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10034_ (.CLK(clknet_leaf_30_mclk),
    .D(_00725_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10035_ (.CLK(clknet_leaf_30_mclk),
    .D(_00726_),
    .RESET_B(net909),
    .Q(\u_glbl_reg.u_random.n1_plus_n0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10036_ (.CLK(clknet_leaf_33_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[19] ),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10037_ (.CLK(clknet_leaf_41_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[20] ),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.n1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10038_ (.CLK(clknet_leaf_34_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[21] ),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.n1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10039_ (.CLK(clknet_leaf_40_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[22] ),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.n1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10040_ (.CLK(clknet_leaf_42_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[23] ),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n1[4] ));
 sky130_fd_sc_hd__dfrtp_2 _10041_ (.CLK(clknet_leaf_36_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[24] ),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.n1[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10042_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[25] ),
    .RESET_B(net950),
    .Q(\u_glbl_reg.u_random.n1[6] ));
 sky130_fd_sc_hd__dfrtp_4 _10043_ (.CLK(clknet_leaf_34_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[26] ),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10044_ (.CLK(clknet_leaf_36_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[27] ),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10045_ (.CLK(clknet_leaf_35_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[28] ),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n1[9] ));
 sky130_fd_sc_hd__dfrtp_2 _10046_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[29] ),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.n1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10047_ (.CLK(clknet_leaf_35_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[30] ),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.n1[11] ));
 sky130_fd_sc_hd__dfrtp_2 _10048_ (.CLK(clknet_leaf_38_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[31] ),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n1[12] ));
 sky130_fd_sc_hd__dfrtp_2 _10049_ (.CLK(clknet_leaf_35_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[0] ),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.n1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10050_ (.CLK(clknet_leaf_37_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[1] ),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10051_ (.CLK(clknet_leaf_34_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[2] ),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10052_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[3] ),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.n1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10053_ (.CLK(clknet_leaf_43_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[4] ),
    .RESET_B(net945),
    .Q(\u_glbl_reg.u_random.n1[17] ));
 sky130_fd_sc_hd__dfrtp_2 _10054_ (.CLK(clknet_leaf_37_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[5] ),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n1[18] ));
 sky130_fd_sc_hd__dfrtp_2 _10055_ (.CLK(clknet_leaf_41_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[6] ),
    .RESET_B(net945),
    .Q(\u_glbl_reg.u_random.n1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10056_ (.CLK(clknet_leaf_40_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[7] ),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.n1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10057_ (.CLK(clknet_leaf_34_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[8] ),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10058_ (.CLK(clknet_leaf_34_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[9] ),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10059_ (.CLK(clknet_leaf_41_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[10] ),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.n1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10060_ (.CLK(clknet_leaf_36_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[11] ),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.n1[24] ));
 sky130_fd_sc_hd__dfrtp_2 _10061_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[12] ),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.n1[25] ));
 sky130_fd_sc_hd__dfrtp_2 _10062_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[13] ),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.n1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10063_ (.CLK(clknet_leaf_36_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[14] ),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10064_ (.CLK(clknet_leaf_35_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[15] ),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n1[28] ));
 sky130_fd_sc_hd__dfrtp_2 _10065_ (.CLK(clknet_leaf_39_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[16] ),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.n1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10066_ (.CLK(clknet_leaf_36_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[17] ),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.n1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10067_ (.CLK(clknet_leaf_38_mclk),
    .D(\u_glbl_reg.u_random.s1_xor_s0[18] ),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n1[31] ));
 sky130_fd_sc_hd__dfrtp_2 _10068_ (.CLK(clknet_leaf_43_mclk),
    .D(_00023_),
    .RESET_B(net943),
    .Q(\u_glbl_reg.u_random.n0[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10069_ (.CLK(clknet_leaf_40_mclk),
    .D(_00024_),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.n0[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10070_ (.CLK(clknet_leaf_34_mclk),
    .D(_00025_),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n0[2] ));
 sky130_fd_sc_hd__dfrtp_4 _10071_ (.CLK(clknet_leaf_39_mclk),
    .D(_00026_),
    .RESET_B(net950),
    .Q(\u_glbl_reg.u_random.n0[3] ));
 sky130_fd_sc_hd__dfrtp_4 _10072_ (.CLK(clknet_leaf_41_mclk),
    .D(_00027_),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.n0[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10073_ (.CLK(clknet_leaf_37_mclk),
    .D(_00028_),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n0[5] ));
 sky130_fd_sc_hd__dfrtp_4 _10074_ (.CLK(clknet_leaf_37_mclk),
    .D(_00029_),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n0[6] ));
 sky130_fd_sc_hd__dfrtp_4 _10075_ (.CLK(clknet_leaf_39_mclk),
    .D(_00030_),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.n0[7] ));
 sky130_fd_sc_hd__dfrtp_2 _10076_ (.CLK(clknet_leaf_36_mclk),
    .D(_00031_),
    .RESET_B(net941),
    .Q(\u_glbl_reg.u_random.n0[8] ));
 sky130_fd_sc_hd__dfrtp_2 _10077_ (.CLK(clknet_leaf_35_mclk),
    .D(_00000_),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n0[9] ));
 sky130_fd_sc_hd__dfrtp_4 _10078_ (.CLK(clknet_leaf_40_mclk),
    .D(_00011_),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.n0[10] ));
 sky130_fd_sc_hd__dfrtp_4 _10079_ (.CLK(clknet_leaf_42_mclk),
    .D(_00015_),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n0[11] ));
 sky130_fd_sc_hd__dfrtp_4 _10080_ (.CLK(clknet_leaf_39_mclk),
    .D(_00016_),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.n0[12] ));
 sky130_fd_sc_hd__dfrtp_4 _10081_ (.CLK(clknet_leaf_40_mclk),
    .D(_00017_),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.n0[13] ));
 sky130_fd_sc_hd__dfrtp_4 _10082_ (.CLK(clknet_leaf_37_mclk),
    .D(_00018_),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.n0[14] ));
 sky130_fd_sc_hd__dfrtp_2 _10083_ (.CLK(clknet_leaf_35_mclk),
    .D(_00019_),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n0[15] ));
 sky130_fd_sc_hd__dfrtp_4 _10084_ (.CLK(clknet_leaf_40_mclk),
    .D(_00020_),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.n0[16] ));
 sky130_fd_sc_hd__dfrtp_2 _10085_ (.CLK(clknet_leaf_42_mclk),
    .D(_00021_),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.n0[17] ));
 sky130_fd_sc_hd__dfrtp_4 _10086_ (.CLK(clknet_leaf_36_mclk),
    .D(_00022_),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.n0[18] ));
 sky130_fd_sc_hd__dfrtp_4 _10087_ (.CLK(clknet_leaf_40_mclk),
    .D(_00001_),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.n0[19] ));
 sky130_fd_sc_hd__dfrtp_4 _10088_ (.CLK(clknet_leaf_42_mclk),
    .D(_00002_),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.n0[20] ));
 sky130_fd_sc_hd__dfrtp_4 _10089_ (.CLK(clknet_leaf_34_mclk),
    .D(_00003_),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n0[21] ));
 sky130_fd_sc_hd__dfrtp_4 _10090_ (.CLK(clknet_leaf_39_mclk),
    .D(_00004_),
    .RESET_B(net954),
    .Q(\u_glbl_reg.u_random.n0[22] ));
 sky130_fd_sc_hd__dfrtp_4 _10091_ (.CLK(clknet_leaf_37_mclk),
    .D(_00005_),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.n0[23] ));
 sky130_fd_sc_hd__dfrtp_2 _10092_ (.CLK(clknet_leaf_35_mclk),
    .D(_00006_),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.n0[24] ));
 sky130_fd_sc_hd__dfrtp_4 _10093_ (.CLK(clknet_leaf_39_mclk),
    .D(_00007_),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.n0[25] ));
 sky130_fd_sc_hd__dfrtp_4 _10094_ (.CLK(clknet_leaf_34_mclk),
    .D(_00008_),
    .RESET_B(net941),
    .Q(\u_glbl_reg.u_random.n0[26] ));
 sky130_fd_sc_hd__dfrtp_2 _10095_ (.CLK(clknet_leaf_36_mclk),
    .D(_00009_),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.n0[27] ));
 sky130_fd_sc_hd__dfrtp_2 _10096_ (.CLK(clknet_leaf_34_mclk),
    .D(_00010_),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.n0[28] ));
 sky130_fd_sc_hd__dfrtp_4 _10097_ (.CLK(clknet_leaf_37_mclk),
    .D(_00012_),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.n0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10098_ (.CLK(clknet_leaf_35_mclk),
    .D(_00013_),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.n0[30] ));
 sky130_fd_sc_hd__dfrtp_4 _10099_ (.CLK(clknet_leaf_38_mclk),
    .D(_00014_),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.n0[31] ));
 sky130_fd_sc_hd__dfrtp_2 _10100_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1856),
    .RESET_B(net943),
    .Q(\u_glbl_reg.u_random.s1[0] ));
 sky130_fd_sc_hd__dfrtp_2 _10101_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1902),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10102_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1857),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.s1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10103_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1871),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.s1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10104_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1858),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.s1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10105_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1877),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.s1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10106_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1904),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.s1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10107_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1914),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10108_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1870),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.s1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10109_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1867),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.s1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10110_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1885),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10111_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1880),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.s1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10112_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1864),
    .RESET_B(net950),
    .Q(\u_glbl_reg.u_random.s1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10113_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1898),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.s1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10114_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1890),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.s1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10115_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1865),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.s1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10116_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1887),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.s1[16] ));
 sky130_fd_sc_hd__dfrtp_2 _10117_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1827),
    .RESET_B(net945),
    .Q(\u_glbl_reg.u_random.s1[17] ));
 sky130_fd_sc_hd__dfrtp_2 _10118_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1882),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.s1[18] ));
 sky130_fd_sc_hd__dfrtp_2 _10119_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1872),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10120_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1860),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.s1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10121_ (.CLK(clknet_2_1__leaf__04359_),
    .D(net1863),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.s1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10122_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1893),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.s1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10123_ (.CLK(clknet_2_3__leaf__04359_),
    .D(net1859),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.s1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10124_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1876),
    .RESET_B(net941),
    .Q(\u_glbl_reg.u_random.s1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10125_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1891),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.s1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10126_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1888),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.s1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10127_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1873),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.s1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10128_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1854),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.s1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10129_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1886),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.s1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10130_ (.CLK(clknet_2_0__leaf__04359_),
    .D(net1866),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.s1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10131_ (.CLK(clknet_2_2__leaf__04359_),
    .D(net1855),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.s1[31] ));
 sky130_fd_sc_hd__dfstp_2 _10132_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1853),
    .SET_B(net943),
    .Q(\u_glbl_reg.u_random.s0[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10133_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1918),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10134_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1883),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.s0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10135_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1916),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.s0[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10136_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1906),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.s0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10137_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1919),
    .RESET_B(net948),
    .Q(\u_glbl_reg.u_random.s0[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10138_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1926),
    .RESET_B(net942),
    .Q(\u_glbl_reg.u_random.s0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10139_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1939),
    .RESET_B(net952),
    .Q(\u_glbl_reg.u_random.s0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10140_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1889),
    .RESET_B(net941),
    .Q(\u_glbl_reg.u_random.s0[8] ));
 sky130_fd_sc_hd__dfrtp_2 _10141_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1881),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.s0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10142_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1908),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.s0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10143_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1907),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.s0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10144_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1929),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.s0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10145_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1940),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.s0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10146_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1909),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.s0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10147_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1874),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.s0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10148_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1917),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.s0[16] ));
 sky130_fd_sc_hd__dfrtp_2 _10149_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1884),
    .RESET_B(net945),
    .Q(\u_glbl_reg.u_random.s0[17] ));
 sky130_fd_sc_hd__dfrtp_2 _10150_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1931),
    .RESET_B(net950),
    .Q(\u_glbl_reg.u_random.s0[18] ));
 sky130_fd_sc_hd__dfrtp_2 _10151_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1927),
    .RESET_B(net954),
    .Q(\u_glbl_reg.u_random.s0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10152_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1901),
    .RESET_B(net951),
    .Q(\u_glbl_reg.u_random.s0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10153_ (.CLK(clknet_2_1__leaf__04358_),
    .D(net1930),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.s0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10154_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1928),
    .RESET_B(net953),
    .Q(\u_glbl_reg.u_random.s0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10155_ (.CLK(clknet_2_3__leaf__04358_),
    .D(net1905),
    .RESET_B(net944),
    .Q(\u_glbl_reg.u_random.s0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10156_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1892),
    .RESET_B(net939),
    .Q(\u_glbl_reg.u_random.s0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10157_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1932),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.s0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10158_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1915),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.s0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10159_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1894),
    .RESET_B(net940),
    .Q(\u_glbl_reg.u_random.s0[27] ));
 sky130_fd_sc_hd__dfrtp_2 _10160_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1897),
    .RESET_B(net937),
    .Q(\u_glbl_reg.u_random.s0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10161_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1912),
    .RESET_B(net947),
    .Q(\u_glbl_reg.u_random.s0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10162_ (.CLK(clknet_2_0__leaf__04358_),
    .D(net1903),
    .RESET_B(net938),
    .Q(\u_glbl_reg.u_random.s0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10163_ (.CLK(clknet_2_2__leaf__04358_),
    .D(net1913),
    .RESET_B(net949),
    .Q(\u_glbl_reg.u_random.s0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10164_ (.CLK(_04391_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.hware_req ),
    .RESET_B(net792),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10165_ (.CLK(_04390_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.hware_req ),
    .RESET_B(net786),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10166_ (.CLK(_04389_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.hware_req ),
    .RESET_B(net915),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10167_ (.CLK(_04388_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.hware_req ),
    .RESET_B(net902),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10168_ (.CLK(_04384_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10169_ (.CLK(_04383_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10170_ (.CLK(_04381_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.hware_req ),
    .RESET_B(net791),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10171_ (.CLK(_04380_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[28].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10172_ (.CLK(_04379_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[27].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10173_ (.CLK(_04378_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[26].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10174_ (.CLK(_04377_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[25].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10175_ (.CLK(_04376_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.hware_req ),
    .RESET_B(net765),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10176_ (.CLK(_04375_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.hware_req ),
    .RESET_B(net902),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[23].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10177_ (.CLK(_04374_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.hware_req ),
    .RESET_B(net906),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10178_ (.CLK(_04373_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.hware_req ),
    .RESET_B(net910),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10179_ (.CLK(_04372_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.hware_req ),
    .RESET_B(net905),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[20].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10180_ (.CLK(_04370_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.hware_req ),
    .RESET_B(net910),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[19].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10181_ (.CLK(_04369_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.hware_req ),
    .RESET_B(net904),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[18].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10182_ (.CLK(_04368_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.hware_req ),
    .RESET_B(net904),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[17].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10183_ (.CLK(_04367_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.hware_req ),
    .RESET_B(net904),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10184_ (.CLK(_04366_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.hware_req ),
    .RESET_B(net807),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10185_ (.CLK(_04365_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.hware_req ),
    .RESET_B(net801),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10186_ (.CLK(_04364_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.hware_req ),
    .RESET_B(net801),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10187_ (.CLK(_04363_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.hware_req ),
    .RESET_B(net784),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10188_ (.CLK(_04362_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.hware_req ),
    .RESET_B(net792),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10189_ (.CLK(_04361_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.hware_req ),
    .RESET_B(net793),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfstp_2 _10190_ (.CLK(clknet_leaf_126_mclk),
    .D(net1654),
    .SET_B(net738),
    .Q(\u_glbl_reg.u_reg_1.flag ));
 sky130_fd_sc_hd__conb_1 _10190__1654 (.LO(net1654));
 sky130_fd_sc_hd__dfrtp_1 _10191_ (.CLK(clknet_1_1__leaf__04395_),
    .D(_00107_),
    .RESET_B(net745),
    .Q(\u_glbl_reg.cfg_rst_ctrl[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10192_ (.CLK(clknet_1_1__leaf__04395_),
    .D(_00108_),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_rst_ctrl[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10193_ (.CLK(clknet_1_0__leaf__04395_),
    .D(_00109_),
    .RESET_B(net735),
    .Q(\u_glbl_reg.cfg_rst_ctrl[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10194_ (.CLK(clknet_1_0__leaf__04395_),
    .D(_00110_),
    .RESET_B(net735),
    .Q(\u_glbl_reg.cfg_rst_ctrl[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10195_ (.CLK(clknet_1_0__leaf__04395_),
    .D(_00111_),
    .RESET_B(net744),
    .Q(\u_glbl_reg.cfg_rst_ctrl[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10196_ (.CLK(clknet_1_0__leaf__04395_),
    .D(_00112_),
    .RESET_B(net738),
    .Q(\u_glbl_reg.cfg_rst_ctrl[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10197_ (.CLK(clknet_1_1__leaf__04395_),
    .D(_00114_),
    .RESET_B(net745),
    .Q(\u_glbl_reg.cfg_rst_ctrl[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10198_ (.CLK(clknet_1_1__leaf__04395_),
    .D(_00115_),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_rst_ctrl[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10199_ (.CLK(clknet_1_0__leaf__04394_),
    .D(_00098_),
    .RESET_B(net783),
    .Q(\u_glbl_reg.cfg_rst_ctrl[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10200_ (.CLK(clknet_1_0__leaf__04394_),
    .D(_00099_),
    .RESET_B(net783),
    .Q(\u_glbl_reg.cfg_rst_ctrl[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10201_ (.CLK(clknet_1_0__leaf__04394_),
    .D(_00100_),
    .RESET_B(net781),
    .Q(\u_glbl_reg.cfg_rst_ctrl[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10202_ (.CLK(clknet_1_1__leaf__04394_),
    .D(_00101_),
    .RESET_B(net782),
    .Q(\u_glbl_reg.cfg_rst_ctrl[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10203_ (.CLK(clknet_1_0__leaf__04394_),
    .D(_00103_),
    .RESET_B(net781),
    .Q(\u_glbl_reg.cfg_rst_ctrl[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10204_ (.CLK(clknet_1_1__leaf__04394_),
    .D(_00104_),
    .RESET_B(net782),
    .Q(\u_glbl_reg.cfg_rst_ctrl[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10205_ (.CLK(clknet_1_1__leaf__04394_),
    .D(_00105_),
    .RESET_B(net783),
    .Q(\u_glbl_reg.cfg_rst_ctrl[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10206_ (.CLK(clknet_1_1__leaf__04394_),
    .D(_00106_),
    .RESET_B(net782),
    .Q(\u_glbl_reg.cfg_rst_ctrl[23] ));
 sky130_fd_sc_hd__dfrtp_4 _10207_ (.CLK(clknet_1_0__leaf__04393_),
    .D(_00121_),
    .RESET_B(net773),
    .Q(\u_glbl_reg.cfg_rst_ctrl[8] ));
 sky130_fd_sc_hd__dfrtp_4 _10208_ (.CLK(clknet_1_0__leaf__04393_),
    .D(_00122_),
    .RESET_B(net773),
    .Q(\u_glbl_reg.cfg_rst_ctrl[9] ));
 sky130_fd_sc_hd__dfrtp_4 _10209_ (.CLK(clknet_1_1__leaf__04393_),
    .D(_00092_),
    .RESET_B(net782),
    .Q(\u_glbl_reg.cfg_rst_ctrl[10] ));
 sky130_fd_sc_hd__dfrtp_4 _10210_ (.CLK(clknet_1_0__leaf__04393_),
    .D(_00093_),
    .RESET_B(net780),
    .Q(\u_glbl_reg.cfg_rst_ctrl[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10211_ (.CLK(clknet_1_0__leaf__04393_),
    .D(_00094_),
    .RESET_B(net777),
    .Q(\u_glbl_reg.cfg_rst_ctrl[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10212_ (.CLK(clknet_1_1__leaf__04393_),
    .D(_00095_),
    .RESET_B(net787),
    .Q(\u_glbl_reg.cfg_rst_ctrl[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10213_ (.CLK(clknet_1_1__leaf__04393_),
    .D(_00096_),
    .RESET_B(net902),
    .Q(\u_glbl_reg.cfg_rst_ctrl[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10214_ (.CLK(clknet_1_1__leaf__04393_),
    .D(_00097_),
    .RESET_B(net787),
    .Q(\u_glbl_reg.cfg_rst_ctrl[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10215_ (.CLK(clknet_1_1__leaf__04392_),
    .D(_00091_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.cfg_rst_ctrl[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10216_ (.CLK(clknet_1_0__leaf__04392_),
    .D(_00102_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.cfg_rst_ctrl[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10217_ (.CLK(clknet_1_0__leaf__04392_),
    .D(_00113_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.cfg_rst_ctrl[2] ));
 sky130_fd_sc_hd__dfrtp_4 _10218_ (.CLK(clknet_1_0__leaf__04392_),
    .D(_00116_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.cfg_rst_ctrl[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10219_ (.CLK(clknet_1_1__leaf__04392_),
    .D(_00117_),
    .RESET_B(net741),
    .Q(\u_glbl_reg.cfg_rst_ctrl[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10220_ (.CLK(clknet_1_0__leaf__04392_),
    .D(_00118_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.cfg_rst_ctrl[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10221_ (.CLK(clknet_1_1__leaf__04392_),
    .D(_00119_),
    .RESET_B(net741),
    .Q(\u_glbl_reg.cfg_rst_ctrl[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10222_ (.CLK(clknet_1_1__leaf__04392_),
    .D(_00120_),
    .RESET_B(net741),
    .Q(\u_glbl_reg.cfg_rst_ctrl[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10223_ (.CLK(clknet_1_1__leaf__04399_),
    .D(net1425),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_15[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10224_ (.CLK(clknet_1_0__leaf__04399_),
    .D(net1418),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_15[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10225_ (.CLK(clknet_1_1__leaf__04399_),
    .D(net1286),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_15[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10226_ (.CLK(clknet_1_0__leaf__04399_),
    .D(net1644),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_15[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10227_ (.CLK(clknet_1_1__leaf__04399_),
    .D(net1636),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_15[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10228_ (.CLK(clknet_1_0__leaf__04399_),
    .D(net1630),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_15[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10229_ (.CLK(clknet_1_1__leaf__04399_),
    .D(net1621),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_15[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10230_ (.CLK(clknet_1_0__leaf__04399_),
    .D(net1613),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_15[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10231_ (.CLK(clknet_1_1__leaf__04398_),
    .D(net1293),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_15[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10232_ (.CLK(clknet_1_0__leaf__04398_),
    .D(net1572),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_15[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10233_ (.CLK(clknet_1_1__leaf__04398_),
    .D(net1488),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_15[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10234_ (.CLK(clknet_1_0__leaf__04398_),
    .D(net1466),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_15[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10235_ (.CLK(clknet_1_1__leaf__04398_),
    .D(net1457),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_15[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10236_ (.CLK(clknet_1_0__leaf__04398_),
    .D(net1448),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_15[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10237_ (.CLK(clknet_1_1__leaf__04398_),
    .D(net1441),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_15[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10238_ (.CLK(clknet_1_0__leaf__04398_),
    .D(net1433),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_15[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10239_ (.CLK(clknet_1_0__leaf__04397_),
    .D(net1534),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10240_ (.CLK(clknet_1_1__leaf__04397_),
    .D(net1526),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10241_ (.CLK(clknet_1_0__leaf__04397_),
    .D(net1519),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10242_ (.CLK(clknet_1_0__leaf__04397_),
    .D(net1512),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10243_ (.CLK(clknet_1_1__leaf__04397_),
    .D(net1505),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10244_ (.CLK(clknet_1_0__leaf__04397_),
    .D(net1498),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_15[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10245_ (.CLK(clknet_1_1__leaf__04397_),
    .D(net1481),
    .RESET_B(net738),
    .Q(\u_glbl_reg.reg_15[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10246_ (.CLK(clknet_1_1__leaf__04397_),
    .D(net1474),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_15[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10247_ (.CLK(clknet_1_1__leaf__04396_),
    .D(net1606),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_15[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10248_ (.CLK(clknet_1_1__leaf__04396_),
    .D(net1598),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10249_ (.CLK(clknet_1_0__leaf__04396_),
    .D(net1589),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10250_ (.CLK(clknet_1_0__leaf__04396_),
    .D(net1582),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10251_ (.CLK(clknet_1_1__leaf__04396_),
    .D(net1566),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10252_ (.CLK(clknet_1_1__leaf__04396_),
    .D(net1559),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_15[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10253_ (.CLK(clknet_1_0__leaf__04396_),
    .D(net1549),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10254_ (.CLK(clknet_1_0__leaf__04396_),
    .D(net1541),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_15[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10255_ (.CLK(clknet_1_0__leaf__04403_),
    .D(net1535),
    .RESET_B(net1044),
    .Q(\u_glbl_reg.reg_16[24] ));
 sky130_fd_sc_hd__dfstp_1 _10256_ (.CLK(clknet_1_1__leaf__04403_),
    .D(net1527),
    .SET_B(net1050),
    .Q(\u_glbl_reg.reg_16[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10257_ (.CLK(clknet_1_1__leaf__04403_),
    .D(net1520),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_16[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10258_ (.CLK(clknet_1_0__leaf__04403_),
    .D(net1512),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_16[27] ));
 sky130_fd_sc_hd__dfstp_1 _10259_ (.CLK(clknet_1_0__leaf__04403_),
    .D(net1505),
    .SET_B(net1048),
    .Q(\u_glbl_reg.reg_16[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10260_ (.CLK(clknet_1_1__leaf__04403_),
    .D(net1501),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_16[29] ));
 sky130_fd_sc_hd__dfstp_1 _10261_ (.CLK(clknet_1_0__leaf__04403_),
    .D(net1481),
    .SET_B(net1048),
    .Q(\u_glbl_reg.reg_16[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10262_ (.CLK(clknet_1_1__leaf__04403_),
    .D(net1474),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_16[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10263_ (.CLK(clknet_1_1__leaf__04402_),
    .D(net1606),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_16[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10264_ (.CLK(clknet_1_1__leaf__04402_),
    .D(net1598),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_16[17] ));
 sky130_fd_sc_hd__dfstp_1 _10265_ (.CLK(clknet_1_1__leaf__04402_),
    .D(net1586),
    .SET_B(net1062),
    .Q(\u_glbl_reg.reg_16[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10266_ (.CLK(clknet_1_1__leaf__04402_),
    .D(net1582),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_16[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10267_ (.CLK(clknet_1_0__leaf__04402_),
    .D(net1564),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_16[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10268_ (.CLK(clknet_1_0__leaf__04402_),
    .D(net1556),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_16[21] ));
 sky130_fd_sc_hd__dfstp_1 _10269_ (.CLK(clknet_1_0__leaf__04402_),
    .D(net1549),
    .SET_B(net1062),
    .Q(\u_glbl_reg.reg_16[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10270_ (.CLK(clknet_1_0__leaf__04402_),
    .D(net1541),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_16[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10271_ (.CLK(clknet_1_1__leaf__04401_),
    .D(net1425),
    .RESET_B(net1060),
    .Q(\u_glbl_reg.reg_16[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10272_ (.CLK(clknet_1_0__leaf__04401_),
    .D(net1418),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_16[9] ));
 sky130_fd_sc_hd__dfstp_1 _10273_ (.CLK(clknet_1_1__leaf__04401_),
    .D(net1288),
    .SET_B(net1069),
    .Q(\u_glbl_reg.reg_16[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10274_ (.CLK(clknet_1_0__leaf__04401_),
    .D(net1645),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_16[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10275_ (.CLK(clknet_1_0__leaf__04401_),
    .D(net1638),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_16[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10276_ (.CLK(clknet_1_0__leaf__04401_),
    .D(net1628),
    .RESET_B(net1060),
    .Q(\u_glbl_reg.reg_16[13] ));
 sky130_fd_sc_hd__dfstp_1 _10277_ (.CLK(clknet_1_1__leaf__04401_),
    .D(net1621),
    .SET_B(net1063),
    .Q(\u_glbl_reg.reg_16[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10278_ (.CLK(clknet_1_1__leaf__04401_),
    .D(net1614),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_16[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10279_ (.CLK(clknet_1_0__leaf__04400_),
    .D(net1293),
    .RESET_B(net1053),
    .Q(\u_glbl_reg.reg_16[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10280_ (.CLK(clknet_1_1__leaf__04400_),
    .D(net1572),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_16[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10281_ (.CLK(clknet_1_0__leaf__04400_),
    .D(net1489),
    .RESET_B(net1053),
    .Q(\u_glbl_reg.reg_16[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10282_ (.CLK(clknet_1_1__leaf__04400_),
    .D(net1466),
    .RESET_B(net1054),
    .Q(\u_glbl_reg.reg_16[3] ));
 sky130_fd_sc_hd__dfstp_1 _10283_ (.CLK(clknet_1_1__leaf__04400_),
    .D(net1458),
    .SET_B(net1054),
    .Q(\u_glbl_reg.reg_16[4] ));
 sky130_fd_sc_hd__dfstp_1 _10284_ (.CLK(clknet_1_1__leaf__04400_),
    .D(net1448),
    .SET_B(net1054),
    .Q(\u_glbl_reg.reg_16[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10285_ (.CLK(clknet_1_0__leaf__04400_),
    .D(net1441),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_16[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10286_ (.CLK(clknet_1_0__leaf__04400_),
    .D(net1433),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_16[7] ));
 sky130_fd_sc_hd__dfstp_1 _10287_ (.CLK(clknet_1_0__leaf__04407_),
    .D(net1293),
    .SET_B(net1052),
    .Q(\u_glbl_reg.reg_17[0] ));
 sky130_fd_sc_hd__dfstp_1 _10288_ (.CLK(clknet_1_1__leaf__04407_),
    .D(net1572),
    .SET_B(net1052),
    .Q(\u_glbl_reg.reg_17[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10289_ (.CLK(clknet_1_0__leaf__04407_),
    .D(net1488),
    .RESET_B(net1047),
    .Q(\u_glbl_reg.reg_17[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10290_ (.CLK(clknet_1_1__leaf__04407_),
    .D(net1466),
    .RESET_B(net1054),
    .Q(\u_glbl_reg.reg_17[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10291_ (.CLK(clknet_1_0__leaf__04407_),
    .D(net1457),
    .RESET_B(net1047),
    .Q(\u_glbl_reg.reg_17[4] ));
 sky130_fd_sc_hd__dfstp_1 _10292_ (.CLK(clknet_1_1__leaf__04407_),
    .D(net1448),
    .SET_B(net1054),
    .Q(\u_glbl_reg.reg_17[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10293_ (.CLK(clknet_1_1__leaf__04407_),
    .D(net1441),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_17[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10294_ (.CLK(clknet_1_0__leaf__04407_),
    .D(net1434),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_17[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10295_ (.CLK(clknet_1_0__leaf__04406_),
    .D(net1427),
    .RESET_B(net1055),
    .Q(\u_glbl_reg.reg_17[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10296_ (.CLK(clknet_1_1__leaf__04406_),
    .D(net1418),
    .RESET_B(net1055),
    .Q(\u_glbl_reg.reg_17[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10297_ (.CLK(clknet_1_1__leaf__04406_),
    .D(net1288),
    .RESET_B(net1069),
    .Q(\u_glbl_reg.reg_17[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10298_ (.CLK(clknet_1_0__leaf__04406_),
    .D(net1644),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_17[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10299_ (.CLK(clknet_1_1__leaf__04406_),
    .D(net1636),
    .RESET_B(net1060),
    .Q(\u_glbl_reg.reg_17[12] ));
 sky130_fd_sc_hd__dfstp_1 _10300_ (.CLK(clknet_1_0__leaf__04406_),
    .D(net1630),
    .SET_B(net1056),
    .Q(\u_glbl_reg.reg_17[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10301_ (.CLK(clknet_1_1__leaf__04406_),
    .D(net1621),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_17[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10302_ (.CLK(clknet_1_0__leaf__04406_),
    .D(net1613),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_17[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10303_ (.CLK(clknet_1_0__leaf__04405_),
    .D(net1534),
    .RESET_B(net1044),
    .Q(\u_glbl_reg.reg_17[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10304_ (.CLK(clknet_1_1__leaf__04405_),
    .D(net1527),
    .RESET_B(net1051),
    .Q(\u_glbl_reg.reg_17[25] ));
 sky130_fd_sc_hd__dfstp_1 _10305_ (.CLK(clknet_1_1__leaf__04405_),
    .D(net1520),
    .SET_B(net1050),
    .Q(\u_glbl_reg.reg_17[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10306_ (.CLK(clknet_1_0__leaf__04405_),
    .D(net1513),
    .RESET_B(net1048),
    .Q(\u_glbl_reg.reg_17[27] ));
 sky130_fd_sc_hd__dfstp_1 _10307_ (.CLK(clknet_1_0__leaf__04405_),
    .D(net1506),
    .SET_B(net1044),
    .Q(\u_glbl_reg.reg_17[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10308_ (.CLK(clknet_1_1__leaf__04405_),
    .D(net1501),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_17[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10309_ (.CLK(clknet_1_1__leaf__04405_),
    .D(net1481),
    .RESET_B(net1048),
    .Q(\u_glbl_reg.reg_17[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10310_ (.CLK(clknet_1_0__leaf__04405_),
    .D(net1474),
    .RESET_B(net1049),
    .Q(\u_glbl_reg.reg_17[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10311_ (.CLK(clknet_1_0__leaf__04404_),
    .D(net1603),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_17[16] ));
 sky130_fd_sc_hd__dfstp_1 _10312_ (.CLK(clknet_1_1__leaf__04404_),
    .D(net1598),
    .SET_B(net1063),
    .Q(\u_glbl_reg.reg_17[17] ));
 sky130_fd_sc_hd__dfstp_1 _10313_ (.CLK(clknet_1_1__leaf__04404_),
    .D(net1589),
    .SET_B(net1062),
    .Q(\u_glbl_reg.reg_17[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10314_ (.CLK(clknet_1_0__leaf__04404_),
    .D(net1579),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_17[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10315_ (.CLK(clknet_1_1__leaf__04404_),
    .D(net1566),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_17[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10316_ (.CLK(clknet_1_0__leaf__04404_),
    .D(net1556),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_17[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10317_ (.CLK(clknet_1_0__leaf__04404_),
    .D(net1549),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_17[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10318_ (.CLK(clknet_1_1__leaf__04404_),
    .D(net1545),
    .RESET_B(net1063),
    .Q(\u_glbl_reg.reg_17[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10319_ (.CLK(clknet_1_1__leaf__04411_),
    .D(net1293),
    .RESET_B(net1053),
    .Q(\u_glbl_reg.reg_18[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10320_ (.CLK(clknet_1_1__leaf__04411_),
    .D(net1572),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_18[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10321_ (.CLK(clknet_1_0__leaf__04411_),
    .D(net1488),
    .RESET_B(net1047),
    .Q(\u_glbl_reg.reg_18[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10322_ (.CLK(clknet_1_1__leaf__04411_),
    .D(net1466),
    .RESET_B(net1053),
    .Q(\u_glbl_reg.reg_18[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10323_ (.CLK(clknet_1_0__leaf__04411_),
    .D(net1457),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.reg_18[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10324_ (.CLK(clknet_1_1__leaf__04411_),
    .D(net1448),
    .RESET_B(net1053),
    .Q(\u_glbl_reg.reg_18[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10325_ (.CLK(clknet_1_0__leaf__04411_),
    .D(net1441),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.reg_18[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10326_ (.CLK(clknet_1_0__leaf__04411_),
    .D(net1434),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_18[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10327_ (.CLK(clknet_1_1__leaf__04410_),
    .D(net1603),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_18[16] ));
 sky130_fd_sc_hd__dfstp_1 _10328_ (.CLK(clknet_1_0__leaf__04410_),
    .D(net1595),
    .SET_B(net1057),
    .Q(\u_glbl_reg.reg_18[17] ));
 sky130_fd_sc_hd__dfstp_1 _10329_ (.CLK(clknet_1_1__leaf__04410_),
    .D(net1586),
    .SET_B(net1058),
    .Q(\u_glbl_reg.reg_18[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10330_ (.CLK(clknet_1_1__leaf__04410_),
    .D(net1579),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_18[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10331_ (.CLK(clknet_1_0__leaf__04410_),
    .D(net1564),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_18[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10332_ (.CLK(clknet_1_0__leaf__04410_),
    .D(net1556),
    .RESET_B(net1057),
    .Q(\u_glbl_reg.reg_18[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10333_ (.CLK(clknet_1_1__leaf__04410_),
    .D(net1549),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_18[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10334_ (.CLK(clknet_1_0__leaf__04410_),
    .D(net1541),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_18[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10335_ (.CLK(clknet_1_0__leaf__04409_),
    .D(net1534),
    .RESET_B(net1044),
    .Q(\u_glbl_reg.reg_18[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10336_ (.CLK(clknet_1_1__leaf__04409_),
    .D(net1527),
    .RESET_B(net1049),
    .Q(\u_glbl_reg.reg_18[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10337_ (.CLK(clknet_1_0__leaf__04409_),
    .D(net1519),
    .RESET_B(net1045),
    .Q(\u_glbl_reg.reg_18[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10338_ (.CLK(clknet_1_0__leaf__04409_),
    .D(net1512),
    .RESET_B(net1045),
    .Q(\u_glbl_reg.reg_18[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10339_ (.CLK(clknet_1_1__leaf__04409_),
    .D(net1506),
    .RESET_B(net1045),
    .Q(\u_glbl_reg.reg_18[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10340_ (.CLK(clknet_1_0__leaf__04409_),
    .D(net1498),
    .RESET_B(net1045),
    .Q(\u_glbl_reg.reg_18[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10341_ (.CLK(clknet_1_1__leaf__04409_),
    .D(net1481),
    .RESET_B(net1049),
    .Q(\u_glbl_reg.reg_18[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10342_ (.CLK(clknet_1_1__leaf__04409_),
    .D(net1474),
    .RESET_B(net1049),
    .Q(\u_glbl_reg.reg_18[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10343_ (.CLK(clknet_1_1__leaf__04408_),
    .D(net1425),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_18[8] ));
 sky130_fd_sc_hd__dfstp_1 _10344_ (.CLK(clknet_1_0__leaf__04408_),
    .D(net1419),
    .SET_B(net1055),
    .Q(\u_glbl_reg.reg_18[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10345_ (.CLK(clknet_1_1__leaf__04408_),
    .D(net1288),
    .RESET_B(net1060),
    .Q(\u_glbl_reg.reg_18[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10346_ (.CLK(clknet_1_0__leaf__04408_),
    .D(net1644),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_18[11] ));
 sky130_fd_sc_hd__dfstp_1 _10347_ (.CLK(clknet_1_1__leaf__04408_),
    .D(net1636),
    .SET_B(net1060),
    .Q(\u_glbl_reg.reg_18[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10348_ (.CLK(clknet_1_0__leaf__04408_),
    .D(net1630),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_18[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10349_ (.CLK(clknet_1_1__leaf__04408_),
    .D(net1621),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_18[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10350_ (.CLK(clknet_1_0__leaf__04408_),
    .D(net1613),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_18[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10351_ (.CLK(clknet_1_1__leaf__04415_),
    .D(net1425),
    .RESET_B(net787),
    .Q(\u_glbl_reg.reg_19[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10352_ (.CLK(clknet_1_0__leaf__04415_),
    .D(net1418),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_19[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10353_ (.CLK(clknet_1_0__leaf__04415_),
    .D(net1286),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_19[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10354_ (.CLK(clknet_1_1__leaf__04415_),
    .D(net1645),
    .RESET_B(net782),
    .Q(\u_glbl_reg.reg_19[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10355_ (.CLK(clknet_1_0__leaf__04415_),
    .D(net1636),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_19[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10356_ (.CLK(clknet_1_1__leaf__04415_),
    .D(net1628),
    .RESET_B(net787),
    .Q(\u_glbl_reg.reg_19[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10357_ (.CLK(clknet_1_0__leaf__04415_),
    .D(net1623),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_19[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10358_ (.CLK(clknet_1_1__leaf__04415_),
    .D(net1615),
    .RESET_B(net787),
    .Q(\u_glbl_reg.reg_19[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10359_ (.CLK(clknet_1_0__leaf__04414_),
    .D(net1293),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_19[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10360_ (.CLK(clknet_1_1__leaf__04414_),
    .D(net1573),
    .RESET_B(net765),
    .Q(\u_glbl_reg.reg_19[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10361_ (.CLK(clknet_1_0__leaf__04414_),
    .D(net1488),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_19[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10362_ (.CLK(clknet_1_1__leaf__04414_),
    .D(net1466),
    .RESET_B(net749),
    .Q(\u_glbl_reg.reg_19[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10363_ (.CLK(clknet_1_0__leaf__04414_),
    .D(net1457),
    .RESET_B(net754),
    .Q(\u_glbl_reg.reg_19[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10364_ (.CLK(clknet_1_0__leaf__04414_),
    .D(net1448),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_19[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10365_ (.CLK(clknet_1_1__leaf__04414_),
    .D(net1442),
    .RESET_B(net750),
    .Q(\u_glbl_reg.reg_19[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10366_ (.CLK(clknet_1_1__leaf__04414_),
    .D(net1434),
    .RESET_B(net750),
    .Q(\u_glbl_reg.reg_19[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10367_ (.CLK(clknet_1_0__leaf__04413_),
    .D(net1535),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_19[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10368_ (.CLK(clknet_1_0__leaf__04413_),
    .D(net1527),
    .RESET_B(net749),
    .Q(\u_glbl_reg.reg_19[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10369_ (.CLK(clknet_1_1__leaf__04413_),
    .D(net1520),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_19[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10370_ (.CLK(clknet_1_1__leaf__04413_),
    .D(net1513),
    .RESET_B(net749),
    .Q(\u_glbl_reg.reg_19[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10371_ (.CLK(clknet_1_0__leaf__04413_),
    .D(net1506),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_19[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10372_ (.CLK(clknet_1_1__leaf__04413_),
    .D(net1501),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_19[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10373_ (.CLK(clknet_1_1__leaf__04413_),
    .D(net1482),
    .RESET_B(net749),
    .Q(\u_glbl_reg.reg_19[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10374_ (.CLK(clknet_1_0__leaf__04413_),
    .D(net1475),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_19[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10375_ (.CLK(clknet_1_0__leaf__04412_),
    .D(net1603),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_19[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10376_ (.CLK(clknet_1_1__leaf__04412_),
    .D(net1598),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_19[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10377_ (.CLK(clknet_1_1__leaf__04412_),
    .D(net1589),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_19[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10378_ (.CLK(clknet_1_0__leaf__04412_),
    .D(net1579),
    .RESET_B(net902),
    .Q(\u_glbl_reg.reg_19[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10379_ (.CLK(clknet_1_1__leaf__04412_),
    .D(net1566),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_19[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10380_ (.CLK(clknet_1_0__leaf__04412_),
    .D(net1556),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_19[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10381_ (.CLK(clknet_1_0__leaf__04412_),
    .D(net1549),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_19[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10382_ (.CLK(clknet_1_1__leaf__04412_),
    .D(net1545),
    .RESET_B(net905),
    .Q(\u_glbl_reg.reg_19[23] ));
 sky130_fd_sc_hd__dfxtp_4 _10383_ (.CLK(clknet_1_1__leaf__04418_),
    .D(_00742_),
    .Q(\u_glbl_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfxtp_2 _10384_ (.CLK(clknet_1_1__leaf__04418_),
    .D(_00743_),
    .Q(\u_glbl_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfxtp_2 _10385_ (.CLK(clknet_1_1__leaf__04418_),
    .D(_00744_),
    .Q(\u_glbl_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfxtp_2 _10386_ (.CLK(clknet_1_1__leaf__04418_),
    .D(_00745_),
    .Q(\u_glbl_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfxtp_1 _10387_ (.CLK(clknet_1_1__leaf__04417_),
    .D(_00746_),
    .Q(\u_glbl_reg.cfg_gpio_dgmode ));
 sky130_fd_sc_hd__dfxtp_1 _10388_ (.CLK(clknet_1_0__leaf__04417_),
    .D(_00747_),
    .Q(\u_glbl_reg.reg_2[9] ));
 sky130_fd_sc_hd__dfxtp_1 _10389_ (.CLK(clknet_1_0__leaf__04417_),
    .D(_00748_),
    .Q(\u_glbl_reg.reg_2[10] ));
 sky130_fd_sc_hd__dfxtp_1 _10390_ (.CLK(clknet_1_1__leaf__04417_),
    .D(_00749_),
    .Q(\u_glbl_reg.reg_2[11] ));
 sky130_fd_sc_hd__dfxtp_1 _10391_ (.CLK(clknet_1_0__leaf__04417_),
    .D(_00750_),
    .Q(\u_glbl_reg.reg_2[12] ));
 sky130_fd_sc_hd__dfxtp_1 _10392_ (.CLK(clknet_1_1__leaf__04417_),
    .D(_00751_),
    .Q(\u_glbl_reg.reg_2[13] ));
 sky130_fd_sc_hd__dfxtp_1 _10393_ (.CLK(clknet_1_0__leaf__04417_),
    .D(_00752_),
    .Q(\u_glbl_reg.reg_2[14] ));
 sky130_fd_sc_hd__dfxtp_1 _10394_ (.CLK(clknet_1_1__leaf__04417_),
    .D(_00753_),
    .Q(\u_glbl_reg.reg_2[15] ));
 sky130_fd_sc_hd__dfxtp_1 _10395_ (.CLK(clknet_1_0__leaf__04416_),
    .D(_00754_),
    .Q(\u_glbl_reg.reg_2[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10396_ (.CLK(clknet_1_0__leaf__04416_),
    .D(_00755_),
    .Q(\u_glbl_reg.reg_2[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10397_ (.CLK(clknet_1_0__leaf__04416_),
    .D(_00756_),
    .Q(\u_glbl_reg.reg_2[2] ));
 sky130_fd_sc_hd__dfxtp_2 _10398_ (.CLK(clknet_1_1__leaf__04416_),
    .D(_00757_),
    .Q(net459));
 sky130_fd_sc_hd__dfxtp_2 _10399_ (.CLK(clknet_1_1__leaf__04416_),
    .D(_00758_),
    .Q(\u_glbl_reg.cfg_mon_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _10400_ (.CLK(clknet_1_1__leaf__04416_),
    .D(_00759_),
    .Q(\u_glbl_reg.cfg_mon_sel[1] ));
 sky130_fd_sc_hd__dfxtp_1 _10401_ (.CLK(clknet_1_1__leaf__04416_),
    .D(_00760_),
    .Q(\u_glbl_reg.cfg_mon_sel[2] ));
 sky130_fd_sc_hd__dfxtp_1 _10402_ (.CLK(clknet_1_0__leaf__04416_),
    .D(_00761_),
    .Q(\u_glbl_reg.cfg_mon_sel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10403_ (.CLK(clknet_1_1__leaf__04423_),
    .D(net1425),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_20[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10404_ (.CLK(clknet_1_0__leaf__04423_),
    .D(net1418),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_20[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10405_ (.CLK(clknet_1_0__leaf__04423_),
    .D(net1288),
    .RESET_B(net788),
    .Q(\u_glbl_reg.reg_20[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10406_ (.CLK(clknet_1_1__leaf__04423_),
    .D(net1645),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_20[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10407_ (.CLK(clknet_1_0__leaf__04423_),
    .D(net1636),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_20[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10408_ (.CLK(clknet_1_1__leaf__04423_),
    .D(net1628),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_20[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10409_ (.CLK(clknet_1_0__leaf__04423_),
    .D(net1623),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_20[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10410_ (.CLK(clknet_1_1__leaf__04423_),
    .D(net1614),
    .RESET_B(net787),
    .Q(\u_glbl_reg.reg_20[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10411_ (.CLK(clknet_1_0__leaf__04422_),
    .D(net1294),
    .RESET_B(net771),
    .Q(\u_glbl_reg.reg_20[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10412_ (.CLK(clknet_1_1__leaf__04422_),
    .D(net1575),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_20[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10413_ (.CLK(clknet_1_0__leaf__04422_),
    .D(net1488),
    .RESET_B(net754),
    .Q(\u_glbl_reg.reg_20[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10414_ (.CLK(clknet_1_1__leaf__04422_),
    .D(net1469),
    .RESET_B(net791),
    .Q(\u_glbl_reg.reg_20[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10415_ (.CLK(clknet_1_0__leaf__04422_),
    .D(net1457),
    .RESET_B(net764),
    .Q(\u_glbl_reg.reg_20[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10416_ (.CLK(clknet_1_1__leaf__04422_),
    .D(net1449),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_20[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10417_ (.CLK(clknet_1_1__leaf__04422_),
    .D(net1442),
    .RESET_B(net794),
    .Q(\u_glbl_reg.reg_20[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10418_ (.CLK(clknet_1_0__leaf__04422_),
    .D(net1433),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_20[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10419_ (.CLK(clknet_1_1__leaf__04421_),
    .D(net1534),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_20[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10420_ (.CLK(clknet_1_1__leaf__04421_),
    .D(net1526),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_20[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10421_ (.CLK(clknet_1_0__leaf__04421_),
    .D(net1519),
    .RESET_B(net741),
    .Q(\u_glbl_reg.reg_20[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10422_ (.CLK(clknet_1_1__leaf__04421_),
    .D(net1512),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_20[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10423_ (.CLK(clknet_1_0__leaf__04421_),
    .D(net1505),
    .RESET_B(net741),
    .Q(\u_glbl_reg.reg_20[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10424_ (.CLK(clknet_1_0__leaf__04421_),
    .D(net1498),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_20[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10425_ (.CLK(clknet_1_0__leaf__04421_),
    .D(net1481),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_20[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10426_ (.CLK(clknet_1_1__leaf__04421_),
    .D(net1474),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_20[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10427_ (.CLK(clknet_1_1__leaf__04420_),
    .D(net1606),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_20[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10428_ (.CLK(clknet_1_1__leaf__04420_),
    .D(net1598),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_20[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10429_ (.CLK(clknet_1_0__leaf__04420_),
    .D(net1589),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_20[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10430_ (.CLK(clknet_1_1__leaf__04420_),
    .D(net1582),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_20[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10431_ (.CLK(clknet_1_1__leaf__04420_),
    .D(net1566),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_20[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10432_ (.CLK(clknet_1_0__leaf__04420_),
    .D(net1556),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_20[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10433_ (.CLK(clknet_1_0__leaf__04420_),
    .D(net1550),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_20[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10434_ (.CLK(clknet_1_0__leaf__04420_),
    .D(net1545),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_20[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10435_ (.CLK(clknet_1_1__leaf__04427_),
    .D(net1425),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_21[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10436_ (.CLK(clknet_1_0__leaf__04427_),
    .D(net1418),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_21[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10437_ (.CLK(clknet_1_0__leaf__04427_),
    .D(net1288),
    .RESET_B(net788),
    .Q(\u_glbl_reg.reg_21[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10438_ (.CLK(clknet_1_1__leaf__04427_),
    .D(net1645),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_21[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10439_ (.CLK(clknet_1_1__leaf__04427_),
    .D(net1636),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_21[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10440_ (.CLK(clknet_1_0__leaf__04427_),
    .D(net1628),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_21[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10441_ (.CLK(clknet_1_0__leaf__04427_),
    .D(net1623),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_21[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10442_ (.CLK(clknet_1_1__leaf__04427_),
    .D(net1614),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_21[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10443_ (.CLK(clknet_1_0__leaf__04426_),
    .D(net1294),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_21[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10444_ (.CLK(clknet_1_1__leaf__04426_),
    .D(net1575),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_21[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10445_ (.CLK(clknet_1_0__leaf__04426_),
    .D(net1488),
    .RESET_B(net754),
    .Q(\u_glbl_reg.reg_21[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10446_ (.CLK(clknet_1_1__leaf__04426_),
    .D(net1469),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_21[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10447_ (.CLK(clknet_1_0__leaf__04426_),
    .D(net1457),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_21[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10448_ (.CLK(clknet_1_1__leaf__04426_),
    .D(net1449),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_21[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10449_ (.CLK(clknet_1_1__leaf__04426_),
    .D(net1442),
    .RESET_B(net765),
    .Q(\u_glbl_reg.reg_21[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10450_ (.CLK(clknet_1_0__leaf__04426_),
    .D(net1433),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_21[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10451_ (.CLK(clknet_1_0__leaf__04425_),
    .D(net1534),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_21[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10452_ (.CLK(clknet_1_1__leaf__04425_),
    .D(net1526),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_21[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10453_ (.CLK(clknet_1_0__leaf__04425_),
    .D(net1519),
    .RESET_B(net741),
    .Q(\u_glbl_reg.reg_21[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10454_ (.CLK(clknet_1_1__leaf__04425_),
    .D(net1513),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_21[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10455_ (.CLK(clknet_1_0__leaf__04425_),
    .D(net1505),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_21[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10456_ (.CLK(clknet_1_0__leaf__04425_),
    .D(net1498),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_21[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10457_ (.CLK(clknet_1_1__leaf__04425_),
    .D(net1482),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_21[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10458_ (.CLK(clknet_1_1__leaf__04425_),
    .D(net1475),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_21[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10459_ (.CLK(clknet_1_0__leaf__04424_),
    .D(net1603),
    .RESET_B(net901),
    .Q(\u_glbl_reg.reg_21[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10460_ (.CLK(clknet_1_1__leaf__04424_),
    .D(net1598),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_21[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10461_ (.CLK(clknet_1_0__leaf__04424_),
    .D(net1589),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_21[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10462_ (.CLK(clknet_1_1__leaf__04424_),
    .D(net1582),
    .RESET_B(net901),
    .Q(\u_glbl_reg.reg_21[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10463_ (.CLK(clknet_1_1__leaf__04424_),
    .D(net1566),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_21[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10464_ (.CLK(clknet_1_1__leaf__04424_),
    .D(net1559),
    .RESET_B(net899),
    .Q(\u_glbl_reg.reg_21[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10465_ (.CLK(clknet_1_0__leaf__04424_),
    .D(net1550),
    .RESET_B(net901),
    .Q(\u_glbl_reg.reg_21[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10466_ (.CLK(clknet_1_0__leaf__04424_),
    .D(net1541),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_21[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10467_ (.CLK(clknet_1_1__leaf__04431_),
    .D(net1425),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_22[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10468_ (.CLK(clknet_1_0__leaf__04431_),
    .D(net1418),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_22[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10469_ (.CLK(clknet_1_0__leaf__04431_),
    .D(net1286),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_22[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10470_ (.CLK(clknet_1_1__leaf__04431_),
    .D(net1645),
    .RESET_B(net782),
    .Q(\u_glbl_reg.reg_22[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10471_ (.CLK(clknet_1_0__leaf__04431_),
    .D(net1636),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_22[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10472_ (.CLK(clknet_1_1__leaf__04431_),
    .D(net1628),
    .RESET_B(net789),
    .Q(\u_glbl_reg.reg_22[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10473_ (.CLK(clknet_1_0__leaf__04431_),
    .D(net1621),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_22[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10474_ (.CLK(clknet_1_1__leaf__04431_),
    .D(net1615),
    .RESET_B(net782),
    .Q(\u_glbl_reg.reg_22[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10475_ (.CLK(clknet_1_0__leaf__04430_),
    .D(net1294),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_22[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10476_ (.CLK(clknet_1_0__leaf__04430_),
    .D(net1573),
    .RESET_B(net750),
    .Q(\u_glbl_reg.reg_22[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10477_ (.CLK(clknet_1_0__leaf__04430_),
    .D(net1488),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_22[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10478_ (.CLK(clknet_1_1__leaf__04430_),
    .D(net1467),
    .RESET_B(net779),
    .Q(\u_glbl_reg.reg_22[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10479_ (.CLK(clknet_1_0__leaf__04430_),
    .D(net1458),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_22[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10480_ (.CLK(clknet_1_1__leaf__04430_),
    .D(net1449),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_22[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10481_ (.CLK(clknet_1_1__leaf__04430_),
    .D(net1442),
    .RESET_B(net779),
    .Q(\u_glbl_reg.reg_22[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10482_ (.CLK(clknet_1_1__leaf__04430_),
    .D(net1434),
    .RESET_B(net750),
    .Q(\u_glbl_reg.reg_22[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10483_ (.CLK(clknet_1_0__leaf__04429_),
    .D(net1534),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_22[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10484_ (.CLK(clknet_1_0__leaf__04429_),
    .D(net1526),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_22[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10485_ (.CLK(clknet_1_1__leaf__04429_),
    .D(net1520),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_22[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10486_ (.CLK(clknet_1_1__leaf__04429_),
    .D(net1513),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_22[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10487_ (.CLK(clknet_1_0__leaf__04429_),
    .D(net1505),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_22[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10488_ (.CLK(clknet_1_1__leaf__04429_),
    .D(net1501),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_22[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10489_ (.CLK(clknet_1_1__leaf__04429_),
    .D(net1482),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_22[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10490_ (.CLK(clknet_1_0__leaf__04429_),
    .D(net1474),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_22[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10491_ (.CLK(clknet_1_1__leaf__04428_),
    .D(net1606),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_22[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10492_ (.CLK(clknet_1_1__leaf__04428_),
    .D(net1598),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_22[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10493_ (.CLK(clknet_1_1__leaf__04428_),
    .D(net1589),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_22[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10494_ (.CLK(clknet_1_0__leaf__04428_),
    .D(net1582),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_22[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10495_ (.CLK(clknet_1_1__leaf__04428_),
    .D(net1566),
    .RESET_B(net908),
    .Q(\u_glbl_reg.reg_22[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10496_ (.CLK(clknet_1_0__leaf__04428_),
    .D(net1559),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_22[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10497_ (.CLK(clknet_1_0__leaf__04428_),
    .D(net1555),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_22[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10498_ (.CLK(clknet_1_0__leaf__04428_),
    .D(net1545),
    .RESET_B(net907),
    .Q(\u_glbl_reg.reg_22[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10499_ (.CLK(clknet_1_0__leaf__04435_),
    .D(net1427),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_23[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10500_ (.CLK(clknet_1_1__leaf__04435_),
    .D(net1418),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_23[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10501_ (.CLK(clknet_1_1__leaf__04435_),
    .D(net1288),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_23[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10502_ (.CLK(clknet_1_0__leaf__04435_),
    .D(net1644),
    .RESET_B(net774),
    .Q(\u_glbl_reg.reg_23[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10503_ (.CLK(clknet_1_1__leaf__04435_),
    .D(net1638),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_23[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10504_ (.CLK(clknet_1_0__leaf__04435_),
    .D(net1630),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_23[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10505_ (.CLK(clknet_1_1__leaf__04435_),
    .D(net1621),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_23[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10506_ (.CLK(clknet_1_0__leaf__04435_),
    .D(net1613),
    .RESET_B(net773),
    .Q(\u_glbl_reg.reg_23[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10507_ (.CLK(clknet_1_1__leaf__04434_),
    .D(net1294),
    .RESET_B(net748),
    .Q(\u_glbl_reg.reg_23[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10508_ (.CLK(clknet_1_1__leaf__04434_),
    .D(net1572),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_23[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10509_ (.CLK(clknet_1_1__leaf__04434_),
    .D(net1489),
    .RESET_B(net765),
    .Q(\u_glbl_reg.reg_23[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10510_ (.CLK(clknet_1_0__leaf__04434_),
    .D(net1466),
    .RESET_B(net753),
    .Q(\u_glbl_reg.reg_23[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10511_ (.CLK(clknet_1_1__leaf__04434_),
    .D(net1458),
    .RESET_B(net763),
    .Q(\u_glbl_reg.reg_23[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10512_ (.CLK(clknet_1_0__leaf__04434_),
    .D(net1448),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_23[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10513_ (.CLK(clknet_1_0__leaf__04434_),
    .D(net1441),
    .RESET_B(net754),
    .Q(\u_glbl_reg.reg_23[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10514_ (.CLK(clknet_1_0__leaf__04434_),
    .D(net1433),
    .RESET_B(net742),
    .Q(\u_glbl_reg.reg_23[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10515_ (.CLK(clknet_1_1__leaf__04433_),
    .D(net1534),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_23[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10516_ (.CLK(clknet_1_0__leaf__04433_),
    .D(net1526),
    .RESET_B(net741),
    .Q(\u_glbl_reg.reg_23[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10517_ (.CLK(clknet_1_0__leaf__04433_),
    .D(net1519),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_23[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10518_ (.CLK(clknet_1_1__leaf__04433_),
    .D(net1512),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_23[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10519_ (.CLK(clknet_1_1__leaf__04433_),
    .D(net1506),
    .RESET_B(net744),
    .Q(\u_glbl_reg.reg_23[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10520_ (.CLK(clknet_1_0__leaf__04433_),
    .D(net1498),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_23[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10521_ (.CLK(clknet_1_0__leaf__04433_),
    .D(net1481),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_23[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10522_ (.CLK(clknet_1_1__leaf__04433_),
    .D(net1475),
    .RESET_B(net747),
    .Q(\u_glbl_reg.reg_23[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10523_ (.CLK(clknet_1_1__leaf__04432_),
    .D(net1603),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_23[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10524_ (.CLK(clknet_1_0__leaf__04432_),
    .D(net1595),
    .RESET_B(net781),
    .Q(\u_glbl_reg.reg_23[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10525_ (.CLK(clknet_1_0__leaf__04432_),
    .D(net1586),
    .RESET_B(net781),
    .Q(\u_glbl_reg.reg_23[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10526_ (.CLK(clknet_1_1__leaf__04432_),
    .D(net1579),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_23[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10527_ (.CLK(clknet_1_0__leaf__04432_),
    .D(net1564),
    .RESET_B(net781),
    .Q(\u_glbl_reg.reg_23[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10528_ (.CLK(clknet_1_0__leaf__04432_),
    .D(net1556),
    .RESET_B(net781),
    .Q(\u_glbl_reg.reg_23[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10529_ (.CLK(clknet_1_1__leaf__04432_),
    .D(net1549),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_23[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10530_ (.CLK(clknet_1_1__leaf__04432_),
    .D(net1541),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_23[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10531_ (.CLK(clknet_1_1__leaf__04439_),
    .D(net1427),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10532_ (.CLK(clknet_1_0__leaf__04439_),
    .D(net1419),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10533_ (.CLK(clknet_1_1__leaf__04439_),
    .D(net1286),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_3[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10534_ (.CLK(clknet_1_1__leaf__04439_),
    .D(net1644),
    .RESET_B(net777),
    .Q(\u_glbl_reg.reg_3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10535_ (.CLK(clknet_1_0__leaf__04439_),
    .D(net1638),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10536_ (.CLK(clknet_1_0__leaf__04439_),
    .D(net1630),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10537_ (.CLK(clknet_1_1__leaf__04439_),
    .D(net1623),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_3[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10538_ (.CLK(clknet_1_0__leaf__04439_),
    .D(net1613),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10539_ (.CLK(clknet_1_1__leaf__04438_),
    .D(net1298),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_3[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10540_ (.CLK(clknet_1_0__leaf__04438_),
    .D(net1575),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10541_ (.CLK(clknet_1_1__leaf__04438_),
    .D(net1496),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_3[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10542_ (.CLK(clknet_1_1__leaf__04438_),
    .D(net1469),
    .RESET_B(net791),
    .Q(\u_glbl_reg.reg_3[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10543_ (.CLK(clknet_1_0__leaf__04438_),
    .D(net1458),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10544_ (.CLK(clknet_1_1__leaf__04438_),
    .D(net1449),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_3[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10545_ (.CLK(clknet_1_0__leaf__04438_),
    .D(net1442),
    .RESET_B(net776),
    .Q(\u_glbl_reg.reg_3[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10546_ (.CLK(clknet_1_0__leaf__04438_),
    .D(net1434),
    .RESET_B(net790),
    .Q(\u_glbl_reg.reg_3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10547_ (.CLK(clknet_1_1__leaf__04437_),
    .D(net1535),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_3[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10548_ (.CLK(clknet_1_0__leaf__04437_),
    .D(net1527),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_3[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10549_ (.CLK(clknet_1_1__leaf__04437_),
    .D(net1520),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_3[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10550_ (.CLK(clknet_1_0__leaf__04437_),
    .D(net1513),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_3[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10551_ (.CLK(clknet_1_0__leaf__04437_),
    .D(net1506),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_3[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10552_ (.CLK(clknet_1_1__leaf__04437_),
    .D(net1499),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_3[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10553_ (.CLK(clknet_1_0__leaf__04437_),
    .D(net1482),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_3[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10554_ (.CLK(clknet_1_1__leaf__04437_),
    .D(net1475),
    .RESET_B(net775),
    .Q(\u_glbl_reg.reg_3[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10555_ (.CLK(clknet_1_0__leaf__04436_),
    .D(net1603),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_3[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10556_ (.CLK(clknet_1_1__leaf__04436_),
    .D(net1598),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_3[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10557_ (.CLK(clknet_1_1__leaf__04436_),
    .D(net1586),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_3[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10558_ (.CLK(clknet_1_1__leaf__04436_),
    .D(net1582),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_3[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10559_ (.CLK(clknet_1_0__leaf__04436_),
    .D(net1564),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_3[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10560_ (.CLK(clknet_1_1__leaf__04436_),
    .D(net1556),
    .RESET_B(net900),
    .Q(\u_glbl_reg.reg_3[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10561_ (.CLK(clknet_1_0__leaf__04436_),
    .D(net1550),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_3[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10562_ (.CLK(clknet_1_0__leaf__04436_),
    .D(net1541),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_3[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10563_ (.CLK(clknet_1_1__leaf__04443_),
    .D(net1534),
    .RESET_B(net746),
    .Q(\u_glbl_reg.cfg_multi_func_sel[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10564_ (.CLK(clknet_1_1__leaf__04443_),
    .D(net1526),
    .RESET_B(net744),
    .Q(\u_glbl_reg.cfg_multi_func_sel[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10565_ (.CLK(clknet_1_0__leaf__04443_),
    .D(net1519),
    .RESET_B(net741),
    .Q(\u_glbl_reg.cfg_multi_func_sel[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10566_ (.CLK(clknet_1_1__leaf__04443_),
    .D(net1512),
    .RESET_B(net747),
    .Q(\u_glbl_reg.cfg_multi_func_sel[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10567_ (.CLK(clknet_1_0__leaf__04443_),
    .D(net1505),
    .RESET_B(net741),
    .Q(\u_glbl_reg.cfg_multi_func_sel[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10568_ (.CLK(clknet_1_0__leaf__04443_),
    .D(net1498),
    .RESET_B(net736),
    .Q(\u_glbl_reg.cfg_multi_func_sel[29] ));
 sky130_fd_sc_hd__dfstp_4 _10569_ (.CLK(clknet_1_1__leaf__04443_),
    .D(net1482),
    .SET_B(net747),
    .Q(\u_glbl_reg.cfg_multi_func_sel[30] ));
 sky130_fd_sc_hd__dfstp_4 _10570_ (.CLK(clknet_1_0__leaf__04443_),
    .D(net1474),
    .SET_B(net741),
    .Q(\u_glbl_reg.cfg_multi_func_sel[31] ));
 sky130_fd_sc_hd__dfrtp_4 _10571_ (.CLK(clknet_1_1__leaf__04442_),
    .D(net1606),
    .RESET_B(net899),
    .Q(\u_glbl_reg.cfg_multi_func_sel[16] ));
 sky130_fd_sc_hd__dfrtp_4 _10572_ (.CLK(clknet_1_1__leaf__04442_),
    .D(net1598),
    .RESET_B(net903),
    .Q(\u_glbl_reg.cfg_multi_func_sel[17] ));
 sky130_fd_sc_hd__dfrtp_4 _10573_ (.CLK(clknet_1_0__leaf__04442_),
    .D(net1586),
    .RESET_B(net902),
    .Q(\u_glbl_reg.cfg_multi_func_sel[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10574_ (.CLK(clknet_1_0__leaf__04442_),
    .D(net1579),
    .RESET_B(net902),
    .Q(\u_glbl_reg.cfg_multi_func_sel[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10575_ (.CLK(clknet_1_1__leaf__04442_),
    .D(net1566),
    .RESET_B(net901),
    .Q(\u_glbl_reg.cfg_multi_func_sel[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10576_ (.CLK(clknet_1_1__leaf__04442_),
    .D(net1559),
    .RESET_B(net903),
    .Q(\u_glbl_reg.cfg_multi_func_sel[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10577_ (.CLK(clknet_1_0__leaf__04442_),
    .D(net1550),
    .RESET_B(net901),
    .Q(\u_glbl_reg.cfg_multi_func_sel[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10578_ (.CLK(clknet_1_0__leaf__04442_),
    .D(net1545),
    .RESET_B(net899),
    .Q(\u_glbl_reg.cfg_multi_func_sel[23] ));
 sky130_fd_sc_hd__dfrtp_4 _10579_ (.CLK(clknet_1_0__leaf__04441_),
    .D(net1427),
    .RESET_B(net777),
    .Q(\u_glbl_reg.cfg_multi_func_sel[8] ));
 sky130_fd_sc_hd__dfrtp_4 _10580_ (.CLK(clknet_1_1__leaf__04441_),
    .D(net1419),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[9] ));
 sky130_fd_sc_hd__dfrtp_4 _10581_ (.CLK(clknet_1_0__leaf__04441_),
    .D(net1286),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10582_ (.CLK(clknet_1_1__leaf__04441_),
    .D(net1643),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10583_ (.CLK(clknet_1_1__leaf__04441_),
    .D(net1638),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[12] ));
 sky130_fd_sc_hd__dfrtp_2 _10584_ (.CLK(clknet_1_0__leaf__04441_),
    .D(net1630),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[13] ));
 sky130_fd_sc_hd__dfrtp_2 _10585_ (.CLK(clknet_1_0__leaf__04441_),
    .D(net1623),
    .RESET_B(net792),
    .Q(\u_glbl_reg.cfg_multi_func_sel[14] ));
 sky130_fd_sc_hd__dfrtp_4 _10586_ (.CLK(clknet_1_1__leaf__04441_),
    .D(net1613),
    .RESET_B(net778),
    .Q(\u_glbl_reg.cfg_multi_func_sel[15] ));
 sky130_fd_sc_hd__dfrtp_4 _10587_ (.CLK(clknet_1_0__leaf__04440_),
    .D(net1294),
    .RESET_B(net764),
    .Q(\u_glbl_reg.cfg_multi_func_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10588_ (.CLK(clknet_1_1__leaf__04440_),
    .D(net1573),
    .RESET_B(net791),
    .Q(\u_glbl_reg.cfg_multi_func_sel[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10589_ (.CLK(clknet_1_0__leaf__04440_),
    .D(net1496),
    .RESET_B(net764),
    .Q(\u_glbl_reg.cfg_multi_func_sel[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10590_ (.CLK(clknet_1_1__leaf__04440_),
    .D(net1467),
    .RESET_B(net794),
    .Q(\u_glbl_reg.cfg_multi_func_sel[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10591_ (.CLK(clknet_1_0__leaf__04440_),
    .D(net1458),
    .RESET_B(net764),
    .Q(\u_glbl_reg.cfg_multi_func_sel[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10592_ (.CLK(clknet_1_1__leaf__04440_),
    .D(net1452),
    .RESET_B(net794),
    .Q(\u_glbl_reg.cfg_multi_func_sel[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10593_ (.CLK(clknet_1_1__leaf__04440_),
    .D(net1442),
    .RESET_B(net791),
    .Q(\u_glbl_reg.cfg_multi_func_sel[6] ));
 sky130_fd_sc_hd__dfrtp_2 _10594_ (.CLK(clknet_1_0__leaf__04440_),
    .D(net1434),
    .RESET_B(net764),
    .Q(\u_glbl_reg.cfg_multi_func_sel[7] ));
 sky130_fd_sc_hd__dfrtp_4 _10595_ (.CLK(clknet_1_1__leaf__04447_),
    .D(net1427),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10596_ (.CLK(clknet_1_1__leaf__04447_),
    .D(net1419),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[1] ));
 sky130_fd_sc_hd__dfrtp_4 _10597_ (.CLK(clknet_1_1__leaf__04447_),
    .D(net1286),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[2] ));
 sky130_fd_sc_hd__dfrtp_4 _10598_ (.CLK(clknet_1_0__leaf__04447_),
    .D(net1644),
    .RESET_B(net750),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[3] ));
 sky130_fd_sc_hd__dfrtp_4 _10599_ (.CLK(clknet_1_0__leaf__04447_),
    .D(net1638),
    .RESET_B(net748),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10600_ (.CLK(clknet_1_1__leaf__04447_),
    .D(net1630),
    .RESET_B(net750),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10601_ (.CLK(clknet_1_0__leaf__04447_),
    .D(net1623),
    .RESET_B(net749),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[6] ));
 sky130_fd_sc_hd__dfrtp_2 _10602_ (.CLK(clknet_1_0__leaf__04447_),
    .D(net1613),
    .RESET_B(net747),
    .Q(\u_glbl_reg.cfg_usb_clk_ctrl[7] ));
 sky130_fd_sc_hd__dfrtp_2 _10603_ (.CLK(clknet_1_0__leaf__04446_),
    .D(net1293),
    .RESET_B(net753),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10604_ (.CLK(clknet_1_1__leaf__04446_),
    .D(net1572),
    .RESET_B(net754),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10605_ (.CLK(clknet_1_1__leaf__04446_),
    .D(net1489),
    .RESET_B(net754),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10606_ (.CLK(clknet_1_1__leaf__04446_),
    .D(net1466),
    .RESET_B(net754),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10607_ (.CLK(clknet_1_1__leaf__04446_),
    .D(net1457),
    .RESET_B(net754),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10608_ (.CLK(clknet_1_0__leaf__04446_),
    .D(net1448),
    .RESET_B(net753),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10609_ (.CLK(clknet_1_0__leaf__04446_),
    .D(net1441),
    .RESET_B(net753),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10610_ (.CLK(clknet_1_0__leaf__04446_),
    .D(net1433),
    .RESET_B(net753),
    .Q(\u_glbl_reg.cfg_rtc_clk_ctrl[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10611_ (.CLK(clknet_1_1__leaf__04445_),
    .D(net1535),
    .RESET_B(net746),
    .Q(\u_glbl_reg.reg_6[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10612_ (.CLK(clknet_1_1__leaf__04445_),
    .D(net1526),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_6[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10613_ (.CLK(clknet_1_0__leaf__04445_),
    .D(net1519),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_6[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10614_ (.CLK(clknet_1_1__leaf__04445_),
    .D(net1513),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_6[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10615_ (.CLK(clknet_1_0__leaf__04445_),
    .D(net1505),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_6[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10616_ (.CLK(clknet_1_0__leaf__04445_),
    .D(net1498),
    .RESET_B(net737),
    .Q(\u_glbl_reg.reg_6[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10617_ (.CLK(clknet_1_0__leaf__04445_),
    .D(net1481),
    .RESET_B(net736),
    .Q(\u_glbl_reg.reg_6[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10618_ (.CLK(clknet_1_1__leaf__04445_),
    .D(net1475),
    .RESET_B(net745),
    .Q(\u_glbl_reg.reg_6[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10619_ (.CLK(clknet_1_0__leaf__04444_),
    .D(net1603),
    .RESET_B(net783),
    .Q(\u_glbl_reg.reg_6[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10620_ (.CLK(clknet_1_0__leaf__04444_),
    .D(net1595),
    .RESET_B(net782),
    .Q(\u_glbl_reg.reg_6[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10621_ (.CLK(clknet_1_1__leaf__04444_),
    .D(net1586),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_6[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10622_ (.CLK(clknet_1_1__leaf__04444_),
    .D(net1579),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_6[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10623_ (.CLK(clknet_1_1__leaf__04444_),
    .D(net1564),
    .RESET_B(net901),
    .Q(\u_glbl_reg.reg_6[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10624_ (.CLK(clknet_1_0__leaf__04444_),
    .D(net1557),
    .RESET_B(net780),
    .Q(\u_glbl_reg.reg_6[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10625_ (.CLK(clknet_1_0__leaf__04444_),
    .D(net1549),
    .RESET_B(net782),
    .Q(\u_glbl_reg.reg_6[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10626_ (.CLK(clknet_1_1__leaf__04444_),
    .D(net1541),
    .RESET_B(net898),
    .Q(\u_glbl_reg.reg_6[23] ));
 sky130_fd_sc_hd__dfrtp_2 _10627_ (.CLK(clknet_1_0__leaf__04451_),
    .D(net1293),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.cfg_ref_pll_div[0] ));
 sky130_fd_sc_hd__dfrtp_4 _10628_ (.CLK(clknet_1_0__leaf__04451_),
    .D(net1572),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.cfg_ref_pll_div[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10629_ (.CLK(clknet_1_0__leaf__04451_),
    .D(net1489),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.cfg_ref_pll_div[2] ));
 sky130_fd_sc_hd__dfstp_2 _10630_ (.CLK(clknet_1_1__leaf__04451_),
    .D(net1467),
    .SET_B(net1054),
    .Q(net226));
 sky130_fd_sc_hd__dfrtp_1 _10631_ (.CLK(clknet_1_1__leaf__04451_),
    .D(net1458),
    .RESET_B(net1054),
    .Q(\u_glbl_reg.reg_7[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10632_ (.CLK(clknet_1_1__leaf__04451_),
    .D(net1449),
    .RESET_B(net1054),
    .Q(\u_glbl_reg.reg_7[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10633_ (.CLK(clknet_1_0__leaf__04451_),
    .D(net1441),
    .RESET_B(net1046),
    .Q(\u_glbl_reg.reg_7[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10634_ (.CLK(clknet_1_1__leaf__04451_),
    .D(net1433),
    .RESET_B(net1052),
    .Q(\u_glbl_reg.reg_7[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10635_ (.CLK(clknet_1_1__leaf__04450_),
    .D(net1535),
    .RESET_B(net1051),
    .Q(\u_glbl_reg.reg_7[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10636_ (.CLK(clknet_1_1__leaf__04450_),
    .D(net1527),
    .RESET_B(net1051),
    .Q(\u_glbl_reg.reg_7[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10637_ (.CLK(clknet_1_0__leaf__04450_),
    .D(net1520),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_7[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10638_ (.CLK(clknet_1_0__leaf__04450_),
    .D(net1513),
    .RESET_B(net1048),
    .Q(\u_glbl_reg.reg_7[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10639_ (.CLK(clknet_1_0__leaf__04450_),
    .D(net1506),
    .RESET_B(net1048),
    .Q(\u_glbl_reg.reg_7[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10640_ (.CLK(clknet_1_1__leaf__04450_),
    .D(net1499),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_7[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10641_ (.CLK(clknet_1_0__leaf__04450_),
    .D(net1482),
    .RESET_B(net1049),
    .Q(\u_glbl_reg.reg_7[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10642_ (.CLK(clknet_1_1__leaf__04450_),
    .D(net1475),
    .RESET_B(net1050),
    .Q(\u_glbl_reg.reg_7[31] ));
 sky130_fd_sc_hd__dfrtp_1 _10643_ (.CLK(clknet_1_0__leaf__04449_),
    .D(net1604),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_7[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10644_ (.CLK(clknet_1_0__leaf__04449_),
    .D(net1595),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_7[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10645_ (.CLK(clknet_1_1__leaf__04449_),
    .D(net1586),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_7[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10646_ (.CLK(clknet_1_0__leaf__04449_),
    .D(net1579),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_7[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10647_ (.CLK(clknet_1_1__leaf__04449_),
    .D(net1564),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_7[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10648_ (.CLK(clknet_1_1__leaf__04449_),
    .D(net1557),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_7[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10649_ (.CLK(clknet_1_0__leaf__04449_),
    .D(net1549),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_7[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10650_ (.CLK(clknet_1_1__leaf__04449_),
    .D(net1541),
    .RESET_B(net1062),
    .Q(\u_glbl_reg.reg_7[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10651_ (.CLK(clknet_1_1__leaf__04448_),
    .D(net1425),
    .RESET_B(net1060),
    .Q(\u_glbl_reg.reg_7[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10652_ (.CLK(clknet_1_0__leaf__04448_),
    .D(net1419),
    .RESET_B(net1057),
    .Q(\u_glbl_reg.reg_7[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10653_ (.CLK(clknet_1_0__leaf__04448_),
    .D(net1286),
    .RESET_B(net1057),
    .Q(\u_glbl_reg.reg_7[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10654_ (.CLK(clknet_1_1__leaf__04448_),
    .D(net1645),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_7[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10655_ (.CLK(clknet_1_0__leaf__04448_),
    .D(net1638),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_7[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10656_ (.CLK(clknet_1_1__leaf__04448_),
    .D(net1628),
    .RESET_B(net1058),
    .Q(\u_glbl_reg.reg_7[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10657_ (.CLK(clknet_1_0__leaf__04448_),
    .D(net1623),
    .RESET_B(net1056),
    .Q(\u_glbl_reg.reg_7[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10658_ (.CLK(clknet_1_1__leaf__04448_),
    .D(net1614),
    .RESET_B(net1059),
    .Q(\u_glbl_reg.reg_7[15] ));
 sky130_fd_sc_hd__dfrtp_4 _10659_ (.CLK(clknet_1_1__leaf__04455_),
    .D(net1540),
    .RESET_B(net1064),
    .Q(net215));
 sky130_fd_sc_hd__dfrtp_4 _10660_ (.CLK(clknet_1_0__leaf__04455_),
    .D(net1532),
    .RESET_B(net1064),
    .Q(net216));
 sky130_fd_sc_hd__dfrtp_4 _10661_ (.CLK(clknet_1_0__leaf__04455_),
    .D(net1525),
    .RESET_B(net1064),
    .Q(net227));
 sky130_fd_sc_hd__dfrtp_4 _10662_ (.CLK(clknet_1_1__leaf__04455_),
    .D(net1518),
    .RESET_B(net1064),
    .Q(net228));
 sky130_fd_sc_hd__dfrtp_4 _10663_ (.CLK(clknet_1_0__leaf__04455_),
    .D(net1511),
    .RESET_B(net1064),
    .Q(net229));
 sky130_fd_sc_hd__dfrtp_4 _10664_ (.CLK(clknet_1_1__leaf__04455_),
    .D(net1504),
    .RESET_B(net1064),
    .Q(net230));
 sky130_fd_sc_hd__dfrtp_4 _10665_ (.CLK(clknet_1_1__leaf__04455_),
    .D(net1487),
    .RESET_B(net1064),
    .Q(net231));
 sky130_fd_sc_hd__dfstp_2 _10666_ (.CLK(clknet_1_0__leaf__04455_),
    .D(net1480),
    .SET_B(net1064),
    .Q(net225));
 sky130_fd_sc_hd__dfrtp_4 _10667_ (.CLK(clknet_1_0__leaf__04454_),
    .D(net1611),
    .RESET_B(net1067),
    .Q(net206));
 sky130_fd_sc_hd__dfrtp_4 _10668_ (.CLK(clknet_1_0__leaf__04454_),
    .D(net1602),
    .RESET_B(net1067),
    .Q(net207));
 sky130_fd_sc_hd__dfrtp_4 _10669_ (.CLK(clknet_1_0__leaf__04454_),
    .D(net1593),
    .RESET_B(net1067),
    .Q(net208));
 sky130_fd_sc_hd__dfrtp_4 _10670_ (.CLK(clknet_1_1__leaf__04454_),
    .D(net1585),
    .RESET_B(net1067),
    .Q(net209));
 sky130_fd_sc_hd__dfrtp_4 _10671_ (.CLK(clknet_1_0__leaf__04454_),
    .D(net1570),
    .RESET_B(net1067),
    .Q(net211));
 sky130_fd_sc_hd__dfrtp_4 _10672_ (.CLK(clknet_1_1__leaf__04454_),
    .D(net1560),
    .RESET_B(net1067),
    .Q(net212));
 sky130_fd_sc_hd__dfrtp_4 _10673_ (.CLK(clknet_1_1__leaf__04454_),
    .D(net1555),
    .RESET_B(net1067),
    .Q(net213));
 sky130_fd_sc_hd__dfrtp_4 _10674_ (.CLK(clknet_1_1__leaf__04454_),
    .D(net1548),
    .RESET_B(net1067),
    .Q(net214));
 sky130_fd_sc_hd__dfstp_4 _10675_ (.CLK(clknet_1_0__leaf__04453_),
    .D(net1429),
    .SET_B(net1066),
    .Q(net223));
 sky130_fd_sc_hd__dfrtp_4 _10676_ (.CLK(clknet_1_1__leaf__04453_),
    .D(net1423),
    .RESET_B(net1066),
    .Q(net224));
 sky130_fd_sc_hd__dfstp_4 _10677_ (.CLK(clknet_1_1__leaf__04453_),
    .D(net1291),
    .SET_B(net1066),
    .Q(net200));
 sky130_fd_sc_hd__dfrtp_4 _10678_ (.CLK(clknet_1_1__leaf__04453_),
    .D(net1647),
    .RESET_B(net1066),
    .Q(net201));
 sky130_fd_sc_hd__dfstp_4 _10679_ (.CLK(clknet_1_1__leaf__04453_),
    .D(net1640),
    .SET_B(net1066),
    .Q(net202));
 sky130_fd_sc_hd__dfrtp_4 _10680_ (.CLK(clknet_1_0__leaf__04453_),
    .D(net1632),
    .RESET_B(net1066),
    .Q(net203));
 sky130_fd_sc_hd__dfrtp_4 _10681_ (.CLK(clknet_1_0__leaf__04453_),
    .D(net1625),
    .RESET_B(net1066),
    .Q(net204));
 sky130_fd_sc_hd__dfrtp_4 _10682_ (.CLK(clknet_1_0__leaf__04453_),
    .D(net1618),
    .RESET_B(net1066),
    .Q(net205));
 sky130_fd_sc_hd__dfstp_2 _10683_ (.CLK(clknet_1_0__leaf__04452_),
    .D(net1302),
    .SET_B(net1065),
    .Q(net199));
 sky130_fd_sc_hd__dfrtp_4 _10684_ (.CLK(clknet_1_0__leaf__04452_),
    .D(net1576),
    .RESET_B(net1065),
    .Q(net210));
 sky130_fd_sc_hd__dfrtp_2 _10685_ (.CLK(clknet_1_1__leaf__04452_),
    .D(net1495),
    .RESET_B(net1065),
    .Q(net217));
 sky130_fd_sc_hd__dfstp_2 _10686_ (.CLK(clknet_1_1__leaf__04452_),
    .D(net1472),
    .SET_B(net1065),
    .Q(net218));
 sky130_fd_sc_hd__dfrtp_4 _10687_ (.CLK(clknet_1_1__leaf__04452_),
    .D(net1462),
    .RESET_B(net1065),
    .Q(net219));
 sky130_fd_sc_hd__dfstp_2 _10688_ (.CLK(clknet_1_0__leaf__04452_),
    .D(net1454),
    .SET_B(net1064),
    .Q(net220));
 sky130_fd_sc_hd__dfstp_2 _10689_ (.CLK(clknet_1_1__leaf__04452_),
    .D(net1446),
    .SET_B(net1064),
    .Q(net221));
 sky130_fd_sc_hd__dfrtp_4 _10690_ (.CLK(clknet_1_0__leaf__04452_),
    .D(net1437),
    .RESET_B(net1065),
    .Q(net222));
 sky130_fd_sc_hd__dfrtp_1 _10691_ (.CLK(\u_glbl_reg.rtc_ref_clk ),
    .D(_00192_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.rtc_clk_div ));
 sky130_fd_sc_hd__dfrtp_1 _10692_ (.CLK(clknet_1_1__leaf__04457_),
    .D(_00195_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.low_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10693_ (.CLK(clknet_1_1__leaf__04457_),
    .D(_00196_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.low_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10694_ (.CLK(clknet_1_0__leaf__04457_),
    .D(_00197_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.low_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10695_ (.CLK(clknet_1_0__leaf__04457_),
    .D(_00198_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.low_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10696_ (.CLK(clknet_1_1__leaf__04457_),
    .D(_00199_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.low_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10697_ (.CLK(clknet_1_0__leaf__04456_),
    .D(_00187_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.high_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10698_ (.CLK(clknet_1_0__leaf__04456_),
    .D(_00188_),
    .RESET_B(net752),
    .Q(\u_glbl_reg.u_rtcclk.high_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10699_ (.CLK(clknet_1_0__leaf__04456_),
    .D(_00189_),
    .RESET_B(net755),
    .Q(\u_glbl_reg.u_rtcclk.high_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10700_ (.CLK(clknet_1_1__leaf__04456_),
    .D(_00190_),
    .RESET_B(net755),
    .Q(\u_glbl_reg.u_rtcclk.high_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10701_ (.CLK(clknet_1_1__leaf__04456_),
    .D(_00191_),
    .RESET_B(net755),
    .Q(\u_glbl_reg.u_rtcclk.high_count[4] ));
 sky130_fd_sc_hd__dlxtn_1 _10702_ (.D(net1306),
    .GATE_N(net1381),
    .Q(\u_glbl_reg.reg_12[0] ));
 sky130_fd_sc_hd__dlxtn_1 _10703_ (.D(net1305),
    .GATE_N(net1381),
    .Q(\u_glbl_reg.reg_12[1] ));
 sky130_fd_sc_hd__dlxtn_1 _10704_ (.D(net1304),
    .GATE_N(net1381),
    .Q(\u_glbl_reg.reg_12[2] ));
 sky130_fd_sc_hd__dlxtn_1 _10705_ (.D(net1650),
    .GATE_N(net1381),
    .Q(\u_glbl_reg.reg_12[3] ));
 sky130_fd_sc_hd__dlxtn_1 _10706_ (.D(net1571),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[4] ));
 sky130_fd_sc_hd__dlxtn_1 _10707_ (.D(net1497),
    .GATE_N(net1383),
    .Q(\u_glbl_reg.reg_12[5] ));
 sky130_fd_sc_hd__dlxtn_1 _10708_ (.D(net1417),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[6] ));
 sky130_fd_sc_hd__dlxtn_1 _10709_ (.D(net1403),
    .GATE_N(net1378),
    .Q(\u_glbl_reg.reg_12[7] ));
 sky130_fd_sc_hd__dlxtn_1 _10710_ (.D(net1397),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[8] ));
 sky130_fd_sc_hd__dlxtn_1 _10711_ (.D(net25),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[9] ));
 sky130_fd_sc_hd__dlxtn_2 _10712_ (.D(net26),
    .GATE_N(net39),
    .Q(\u_glbl_reg.reg_12[10] ));
 sky130_fd_sc_hd__dlxtn_4 _10713_ (.D(net27),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[11] ));
 sky130_fd_sc_hd__dlxtn_2 _10714_ (.D(net1396),
    .GATE_N(net1379),
    .Q(\u_glbl_reg.reg_12[12] ));
 sky130_fd_sc_hd__dlxtn_2 _10715_ (.D(net1394),
    .GATE_N(net1378),
    .Q(\u_glbl_reg.reg_12[13] ));
 sky130_fd_sc_hd__dlxtn_1 _10716_ (.D(net1391),
    .GATE_N(net1378),
    .Q(\u_glbl_reg.reg_12[14] ));
 sky130_fd_sc_hd__dlxtn_1 _10717_ (.D(net1390),
    .GATE_N(net1384),
    .Q(\u_glbl_reg.reg_12[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10718_ (.CLK(_04462_),
    .D(_00224_),
    .RESET_B(net1378),
    .Q(net489));
 sky130_fd_sc_hd__dfrtp_1 _10719_ (.CLK(clknet_1_0__leaf__04461_),
    .D(_00216_),
    .RESET_B(net1378),
    .Q(net481));
 sky130_fd_sc_hd__dfrtp_1 _10720_ (.CLK(clknet_1_1__leaf__04461_),
    .D(_00217_),
    .RESET_B(net1378),
    .Q(net482));
 sky130_fd_sc_hd__dfrtp_1 _10721_ (.CLK(clknet_1_0__leaf__04461_),
    .D(_00218_),
    .RESET_B(net1378),
    .Q(net483));
 sky130_fd_sc_hd__dfrtp_1 _10722_ (.CLK(clknet_1_1__leaf__04461_),
    .D(_00219_),
    .RESET_B(net1379),
    .Q(net484));
 sky130_fd_sc_hd__dfrtp_2 _10723_ (.CLK(clknet_1_0__leaf__04461_),
    .D(_00220_),
    .RESET_B(net1378),
    .Q(net485));
 sky130_fd_sc_hd__dfrtp_1 _10724_ (.CLK(clknet_1_1__leaf__04461_),
    .D(_00221_),
    .RESET_B(net1378),
    .Q(net486));
 sky130_fd_sc_hd__dfrtp_2 _10725_ (.CLK(clknet_1_0__leaf__04461_),
    .D(_00223_),
    .RESET_B(net1378),
    .Q(net488));
 sky130_fd_sc_hd__dfrtp_4 _10726_ (.CLK(clknet_1_1__leaf__04460_),
    .D(_00207_),
    .RESET_B(net1382),
    .Q(net472));
 sky130_fd_sc_hd__dfrtp_1 _10727_ (.CLK(clknet_1_0__leaf__04460_),
    .D(_00208_),
    .RESET_B(net1379),
    .Q(net473));
 sky130_fd_sc_hd__dfrtp_4 _10728_ (.CLK(clknet_1_1__leaf__04460_),
    .D(_00209_),
    .RESET_B(net1382),
    .Q(net474));
 sky130_fd_sc_hd__dfrtp_4 _10729_ (.CLK(clknet_1_0__leaf__04460_),
    .D(_00210_),
    .RESET_B(net1379),
    .Q(net475));
 sky130_fd_sc_hd__dfrtp_4 _10730_ (.CLK(clknet_1_1__leaf__04460_),
    .D(_00212_),
    .RESET_B(net1382),
    .Q(net477));
 sky130_fd_sc_hd__dfrtp_4 _10731_ (.CLK(clknet_1_0__leaf__04460_),
    .D(_00213_),
    .RESET_B(net1379),
    .Q(net478));
 sky130_fd_sc_hd__dfrtp_4 _10732_ (.CLK(clknet_1_0__leaf__04460_),
    .D(_00214_),
    .RESET_B(net1379),
    .Q(net479));
 sky130_fd_sc_hd__dfrtp_4 _10733_ (.CLK(clknet_1_1__leaf__04460_),
    .D(_00215_),
    .RESET_B(net1379),
    .Q(net480));
 sky130_fd_sc_hd__dfrtp_4 _10734_ (.CLK(clknet_1_1__leaf__04459_),
    .D(_00230_),
    .RESET_B(net1382),
    .Q(net495));
 sky130_fd_sc_hd__dfrtp_4 _10735_ (.CLK(clknet_1_0__leaf__04459_),
    .D(_00231_),
    .RESET_B(net1382),
    .Q(net496));
 sky130_fd_sc_hd__dfrtp_4 _10736_ (.CLK(clknet_1_1__leaf__04459_),
    .D(_00201_),
    .RESET_B(net1382),
    .Q(net466));
 sky130_fd_sc_hd__dfrtp_4 _10737_ (.CLK(clknet_1_1__leaf__04459_),
    .D(_00202_),
    .RESET_B(net1382),
    .Q(net467));
 sky130_fd_sc_hd__dfrtp_4 _10738_ (.CLK(clknet_1_0__leaf__04459_),
    .D(_00203_),
    .RESET_B(net1382),
    .Q(net468));
 sky130_fd_sc_hd__dfrtp_4 _10739_ (.CLK(clknet_1_0__leaf__04459_),
    .D(_00204_),
    .RESET_B(net1382),
    .Q(net469));
 sky130_fd_sc_hd__dfrtp_4 _10740_ (.CLK(clknet_1_0__leaf__04459_),
    .D(_00205_),
    .RESET_B(net1382),
    .Q(net470));
 sky130_fd_sc_hd__dfrtp_4 _10741_ (.CLK(clknet_1_1__leaf__04459_),
    .D(_00206_),
    .RESET_B(net1383),
    .Q(net471));
 sky130_fd_sc_hd__dfrtp_2 _10742_ (.CLK(clknet_1_1__leaf__04458_),
    .D(_00200_),
    .RESET_B(net1381),
    .Q(net465));
 sky130_fd_sc_hd__dfrtp_4 _10743_ (.CLK(clknet_1_0__leaf__04458_),
    .D(_00211_),
    .RESET_B(net1380),
    .Q(net476));
 sky130_fd_sc_hd__dfrtp_2 _10744_ (.CLK(clknet_1_1__leaf__04458_),
    .D(_00222_),
    .RESET_B(net1380),
    .Q(net487));
 sky130_fd_sc_hd__dfrtp_4 _10745_ (.CLK(clknet_1_0__leaf__04458_),
    .D(_00225_),
    .RESET_B(net1380),
    .Q(net490));
 sky130_fd_sc_hd__dfrtp_4 _10746_ (.CLK(clknet_1_1__leaf__04458_),
    .D(_00226_),
    .RESET_B(net1381),
    .Q(net491));
 sky130_fd_sc_hd__dfrtp_2 _10747_ (.CLK(clknet_1_0__leaf__04458_),
    .D(_00227_),
    .RESET_B(net1380),
    .Q(net492));
 sky130_fd_sc_hd__dfrtp_4 _10748_ (.CLK(clknet_1_1__leaf__04458_),
    .D(_00228_),
    .RESET_B(net1380),
    .Q(net493));
 sky130_fd_sc_hd__dfrtp_2 _10749_ (.CLK(clknet_1_0__leaf__04458_),
    .D(_00229_),
    .RESET_B(net1380),
    .Q(net494));
 sky130_fd_sc_hd__dfrtp_1 _10750_ (.CLK(\u_glbl_reg.u_usb_clk_sel.A0 ),
    .D(_00242_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usb_clk_sel.A1 ));
 sky130_fd_sc_hd__dfrtp_1 _10751_ (.CLK(clknet_1_1__leaf__04464_),
    .D(_00245_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.u_usbclk.low_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10752_ (.CLK(clknet_1_1__leaf__04464_),
    .D(_00246_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.u_usbclk.low_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10753_ (.CLK(clknet_1_1__leaf__04464_),
    .D(_00247_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.u_usbclk.low_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10754_ (.CLK(clknet_1_0__leaf__04464_),
    .D(_00248_),
    .RESET_B(net739),
    .Q(\u_glbl_reg.u_usbclk.low_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10755_ (.CLK(clknet_1_0__leaf__04464_),
    .D(_00249_),
    .RESET_B(net743),
    .Q(\u_glbl_reg.u_usbclk.low_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10756_ (.CLK(clknet_1_1__leaf__04463_),
    .D(_00237_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usbclk.high_count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10757_ (.CLK(clknet_1_1__leaf__04463_),
    .D(_00238_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usbclk.high_count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10758_ (.CLK(clknet_1_0__leaf__04463_),
    .D(_00239_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usbclk.high_count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10759_ (.CLK(clknet_1_0__leaf__04463_),
    .D(_00240_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usbclk.high_count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10760_ (.CLK(clknet_1_0__leaf__04463_),
    .D(_00241_),
    .RESET_B(net740),
    .Q(\u_glbl_reg.u_usbclk.high_count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10761_ (.CLK(clknet_2_1__leaf__04353_),
    .D(net2318),
    .RESET_B(net915),
    .Q(\u_glbl_reg.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10762_ (.CLK(clknet_2_1__leaf__04353_),
    .D(net2063),
    .RESET_B(net805),
    .Q(\u_glbl_reg.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10763_ (.CLK(clknet_2_1__leaf__04353_),
    .D(\u_glbl_reg.reg_out[2] ),
    .RESET_B(net805),
    .Q(\u_glbl_reg.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10764_ (.CLK(clknet_2_3__leaf__04353_),
    .D(\u_glbl_reg.reg_out[3] ),
    .RESET_B(net916),
    .Q(\u_glbl_reg.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10765_ (.CLK(clknet_2_3__leaf__04353_),
    .D(\u_glbl_reg.reg_out[4] ),
    .RESET_B(net915),
    .Q(\u_glbl_reg.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10766_ (.CLK(clknet_2_1__leaf__04353_),
    .D(\u_glbl_reg.reg_out[5] ),
    .RESET_B(net915),
    .Q(\u_glbl_reg.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10767_ (.CLK(clknet_2_1__leaf__04353_),
    .D(\u_glbl_reg.reg_out[6] ),
    .RESET_B(net801),
    .Q(\u_glbl_reg.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10768_ (.CLK(clknet_2_1__leaf__04353_),
    .D(\u_glbl_reg.reg_out[7] ),
    .RESET_B(net801),
    .Q(\u_glbl_reg.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10769_ (.CLK(clknet_2_3__leaf__04353_),
    .D(net1961),
    .RESET_B(net906),
    .Q(\u_glbl_reg.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10770_ (.CLK(clknet_2_3__leaf__04353_),
    .D(net2033),
    .RESET_B(net902),
    .Q(\u_glbl_reg.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10771_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net2052),
    .RESET_B(net902),
    .Q(\u_glbl_reg.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10772_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net1983),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10773_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net1992),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10774_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net1966),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10775_ (.CLK(clknet_2_3__leaf__04353_),
    .D(net1994),
    .RESET_B(net902),
    .Q(\u_glbl_reg.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10776_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net1969),
    .RESET_B(net786),
    .Q(\u_glbl_reg.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10777_ (.CLK(clknet_2_2__leaf__04353_),
    .D(\u_glbl_reg.reg_out[16] ),
    .RESET_B(net904),
    .Q(\u_glbl_reg.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10778_ (.CLK(clknet_2_2__leaf__04353_),
    .D(\u_glbl_reg.reg_out[17] ),
    .RESET_B(net905),
    .Q(\u_glbl_reg.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10779_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2010),
    .RESET_B(net910),
    .Q(\u_glbl_reg.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10780_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net1986),
    .RESET_B(net910),
    .Q(\u_glbl_reg.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10781_ (.CLK(clknet_2_2__leaf__04353_),
    .D(\u_glbl_reg.reg_out[20] ),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10782_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2057),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10783_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2026),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10784_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net1997),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10785_ (.CLK(clknet_2_3__leaf__04353_),
    .D(net2015),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10786_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net2279),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_2 _10787_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2005),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10788_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2037),
    .RESET_B(net903),
    .Q(\u_glbl_reg.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_2 _10789_ (.CLK(clknet_2_2__leaf__04353_),
    .D(net2020),
    .RESET_B(net912),
    .Q(\u_glbl_reg.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10790_ (.CLK(clknet_2_0__leaf__04353_),
    .D(net2002),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10791_ (.CLK(clknet_2_0__leaf__04353_),
    .D(\u_glbl_reg.reg_out[30] ),
    .RESET_B(net785),
    .Q(\u_glbl_reg.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10792_ (.CLK(clknet_2_0__leaf__04353_),
    .D(\u_glbl_reg.reg_out[31] ),
    .RESET_B(net784),
    .Q(\u_glbl_reg.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_4 _10793_ (.CLK(clknet_leaf_22_mclk),
    .D(_00038_),
    .RESET_B(net929),
    .Q(\u_glbl_reg.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _10794_ (.CLK(clknet_leaf_127_mclk),
    .D(net196),
    .RESET_B(net738),
    .Q(\u_glbl_reg.usb_intr_s ));
 sky130_fd_sc_hd__dfrtp_2 _10795_ (.CLK(clknet_leaf_126_mclk),
    .D(net2198),
    .RESET_B(net739),
    .Q(\u_glbl_reg.usb_intr_ss ));
 sky130_fd_sc_hd__dfrtp_1 _10796_ (.CLK(clknet_leaf_127_mclk),
    .D(net44),
    .RESET_B(net738),
    .Q(\u_glbl_reg.i2cm_intr_s ));
 sky130_fd_sc_hd__dfrtp_2 _10797_ (.CLK(clknet_leaf_126_mclk),
    .D(net2195),
    .RESET_B(net739),
    .Q(\u_glbl_reg.i2cm_intr_ss ));
 sky130_fd_sc_hd__dfrtp_1 _10798_ (.CLK(clknet_leaf_44_mclk),
    .D(net133),
    .RESET_B(net959),
    .Q(\u_glbl_reg.rtc_intr_s ));
 sky130_fd_sc_hd__dfrtp_2 _10799_ (.CLK(clknet_leaf_44_mclk),
    .D(net2313),
    .RESET_B(net957),
    .Q(\u_glbl_reg.rtc_intr_ss ));
 sky130_fd_sc_hd__dfrtp_1 _10800_ (.CLK(clknet_leaf_46_mclk),
    .D(net46),
    .RESET_B(net968),
    .Q(\u_glbl_reg.ir_intr_s ));
 sky130_fd_sc_hd__dfrtp_2 _10801_ (.CLK(clknet_leaf_44_mclk),
    .D(\u_glbl_reg.ir_intr_s ),
    .RESET_B(net957),
    .Q(\u_glbl_reg.ir_intr_ss ));
 sky130_fd_sc_hd__dfrtp_1 _10802_ (.CLK(clknet_1_1__leaf__04550_),
    .D(net1825),
    .RESET_B(net1000),
    .Q(\u_pwm.reg_rdata_glbl[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10803_ (.CLK(clknet_1_1__leaf__04550_),
    .D(net1823),
    .RESET_B(net888),
    .Q(\u_pwm.reg_rdata_glbl[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10804_ (.CLK(clknet_1_1__leaf__04550_),
    .D(net1835),
    .RESET_B(net888),
    .Q(\u_pwm.reg_rdata_glbl[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10805_ (.CLK(clknet_1_1__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[3] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_glbl[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10806_ (.CLK(clknet_1_1__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[4] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_glbl[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10807_ (.CLK(clknet_1_1__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[5] ),
    .RESET_B(net1011),
    .Q(\u_pwm.reg_rdata_glbl[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10808_ (.CLK(clknet_1_1__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[8] ),
    .RESET_B(net999),
    .Q(\u_pwm.reg_rdata_glbl[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10809_ (.CLK(clknet_1_0__leaf__04550_),
    .D(net1817),
    .RESET_B(net877),
    .Q(\u_pwm.reg_rdata_glbl[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10810_ (.CLK(clknet_1_0__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[10] ),
    .RESET_B(net876),
    .Q(\u_pwm.reg_rdata_glbl[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10811_ (.CLK(clknet_1_0__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[16] ),
    .RESET_B(net982),
    .Q(\u_pwm.reg_rdata_glbl[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10812_ (.CLK(clknet_1_0__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[17] ),
    .RESET_B(net875),
    .Q(\u_pwm.reg_rdata_glbl[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10813_ (.CLK(clknet_1_0__leaf__04550_),
    .D(\u_pwm.u_glbl_reg.reg_out[18] ),
    .RESET_B(net981),
    .Q(\u_pwm.reg_rdata_glbl[18] ));
 sky130_fd_sc_hd__dlclkp_1 _10814_ (.CLK(clknet_leaf_56_mclk),
    .GATE(net1307),
    .GCLK(_04347_));
 sky130_fd_sc_hd__dfrtp_2 _10815_ (.CLK(clknet_1_0__leaf__04347_),
    .D(net1342),
    .RESET_B(net924),
    .Q(\reg_blk_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10816_ (.CLK(clknet_1_0__leaf__04347_),
    .D(net1341),
    .RESET_B(net924),
    .Q(\reg_blk_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10817_ (.CLK(clknet_1_1__leaf__04347_),
    .D(net1340),
    .RESET_B(net923),
    .Q(\reg_blk_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10818_ (.CLK(clknet_1_1__leaf__04347_),
    .D(net1374),
    .RESET_B(net924),
    .Q(\reg_blk_sel[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10819_ (.CLK(_04387_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.hware_req ),
    .RESET_B(net804),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10820_ (.CLK(_04386_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.hware_req ),
    .RESET_B(net776),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10821_ (.CLK(_04385_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.hware_req ),
    .RESET_B(net776),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10822_ (.CLK(_04382_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .RESET_B(net915),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_4 _10823_ (.CLK(_04371_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .RESET_B(net902),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_2 _10824_ (.CLK(_04360_),
    .D(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .RESET_B(net915),
    .Q(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10825_ (.CLK(clknet_leaf_63_mclk),
    .D(_00578_),
    .RESET_B(net1018),
    .Q(\u_ws281x.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _10826_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[0] ),
    .RESET_B(net1018),
    .Q(\u_ws281x.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10827_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[1] ),
    .RESET_B(net1018),
    .Q(\u_ws281x.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10828_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[2] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10829_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[3] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _10830_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[4] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10831_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[5] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10832_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[6] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10833_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[7] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10834_ (.CLK(clknet_2_3__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[8] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _10835_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[9] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10836_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[10] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10837_ (.CLK(clknet_2_3__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[11] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10838_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[12] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10839_ (.CLK(clknet_2_3__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[13] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _10840_ (.CLK(clknet_2_3__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[14] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10841_ (.CLK(clknet_2_3__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[15] ),
    .RESET_B(net1024),
    .Q(\u_ws281x.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _10842_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[16] ),
    .RESET_B(net963),
    .Q(\u_ws281x.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _10843_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[17] ),
    .RESET_B(net1020),
    .Q(\u_ws281x.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _10844_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[18] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _10845_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[19] ),
    .RESET_B(net971),
    .Q(\u_ws281x.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _10846_ (.CLK(clknet_2_1__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[20] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _10847_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[21] ),
    .RESET_B(net971),
    .Q(\u_ws281x.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _10848_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[22] ),
    .RESET_B(net1019),
    .Q(\u_ws281x.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _10849_ (.CLK(clknet_2_0__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[23] ),
    .RESET_B(net971),
    .Q(\u_ws281x.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _10850_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[24] ),
    .RESET_B(net1026),
    .Q(\u_ws281x.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _10851_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[25] ),
    .RESET_B(net1026),
    .Q(\u_ws281x.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _10852_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[26] ),
    .RESET_B(net972),
    .Q(\u_ws281x.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _10853_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[27] ),
    .RESET_B(net973),
    .Q(\u_ws281x.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _10854_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[28] ),
    .RESET_B(net1026),
    .Q(\u_ws281x.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _10855_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[29] ),
    .RESET_B(net973),
    .Q(\u_ws281x.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _10856_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[30] ),
    .RESET_B(net973),
    .Q(\u_ws281x.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10857_ (.CLK(clknet_2_2__leaf__04653_),
    .D(\u_ws281x.u_reg.reg_out[31] ),
    .RESET_B(net973),
    .Q(\u_ws281x.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_2 _10858_ (.CLK(clknet_1_1__leaf__04672_),
    .D(net1609),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th0_period[6] ));
 sky130_fd_sc_hd__dfrtp_4 _10859_ (.CLK(clknet_1_0__leaf__04672_),
    .D(net1601),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th0_period[7] ));
 sky130_fd_sc_hd__dfrtp_4 _10860_ (.CLK(clknet_1_0__leaf__04672_),
    .D(net1591),
    .RESET_B(net1024),
    .Q(\u_ws281x.cfg_th0_period[8] ));
 sky130_fd_sc_hd__dfrtp_4 _10861_ (.CLK(clknet_1_0__leaf__04672_),
    .D(net1583),
    .RESET_B(net1024),
    .Q(\u_ws281x.cfg_th0_period[9] ));
 sky130_fd_sc_hd__dfrtp_2 _10862_ (.CLK(clknet_1_0__leaf__04672_),
    .D(net1570),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th1_period[0] ));
 sky130_fd_sc_hd__dfrtp_2 _10863_ (.CLK(clknet_1_1__leaf__04672_),
    .D(net1563),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th1_period[1] ));
 sky130_fd_sc_hd__dfrtp_4 _10864_ (.CLK(clknet_1_1__leaf__04672_),
    .D(net1554),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th1_period[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10865_ (.CLK(clknet_1_1__leaf__04672_),
    .D(net1546),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th1_period[3] ));
 sky130_fd_sc_hd__dfrtp_4 _10866_ (.CLK(clknet_1_1__leaf__04673_),
    .D(net1540),
    .RESET_B(net1026),
    .Q(\u_ws281x.cfg_th1_period[4] ));
 sky130_fd_sc_hd__dfrtp_4 _10867_ (.CLK(clknet_1_0__leaf__04673_),
    .D(net1532),
    .RESET_B(net1026),
    .Q(\u_ws281x.cfg_th1_period[5] ));
 sky130_fd_sc_hd__dfrtp_4 _10868_ (.CLK(clknet_1_0__leaf__04673_),
    .D(net1525),
    .RESET_B(net972),
    .Q(\u_ws281x.cfg_th1_period[6] ));
 sky130_fd_sc_hd__dfrtp_4 _10869_ (.CLK(clknet_1_0__leaf__04673_),
    .D(net1518),
    .RESET_B(net971),
    .Q(\u_ws281x.cfg_th1_period[7] ));
 sky130_fd_sc_hd__dfrtp_4 _10870_ (.CLK(clknet_1_1__leaf__04673_),
    .D(net1511),
    .RESET_B(net1026),
    .Q(\u_ws281x.cfg_th1_period[8] ));
 sky130_fd_sc_hd__dfrtp_4 _10871_ (.CLK(clknet_1_0__leaf__04673_),
    .D(net1504),
    .RESET_B(net973),
    .Q(\u_ws281x.cfg_th1_period[9] ));
 sky130_fd_sc_hd__dfrtp_1 _10872_ (.CLK(clknet_1_1__leaf__04673_),
    .D(net1487),
    .RESET_B(net973),
    .Q(\u_ws281x.u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _10873_ (.CLK(clknet_1_1__leaf__04673_),
    .D(net1480),
    .RESET_B(net973),
    .Q(\u_ws281x.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_2 _10874_ (.CLK(clknet_1_0__leaf__04674_),
    .D(net1302),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_clk_period[0] ));
 sky130_fd_sc_hd__dfrtp_2 _10875_ (.CLK(clknet_1_0__leaf__04674_),
    .D(net1576),
    .RESET_B(net1031),
    .Q(\u_ws281x.cfg_clk_period[1] ));
 sky130_fd_sc_hd__dfrtp_1 _10876_ (.CLK(clknet_1_0__leaf__04674_),
    .D(net1493),
    .RESET_B(net1031),
    .Q(\u_ws281x.cfg_clk_period[2] ));
 sky130_fd_sc_hd__dfrtp_1 _10877_ (.CLK(clknet_1_0__leaf__04674_),
    .D(net1470),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_clk_period[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10878_ (.CLK(clknet_1_1__leaf__04674_),
    .D(net1462),
    .RESET_B(net1022),
    .Q(\u_ws281x.cfg_clk_period[4] ));
 sky130_fd_sc_hd__dfrtp_2 _10879_ (.CLK(clknet_1_1__leaf__04674_),
    .D(net1453),
    .RESET_B(net1034),
    .Q(\u_ws281x.cfg_clk_period[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10880_ (.CLK(clknet_1_1__leaf__04674_),
    .D(net1446),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_clk_period[6] ));
 sky130_fd_sc_hd__dfrtp_2 _10881_ (.CLK(clknet_1_1__leaf__04674_),
    .D(net1437),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_clk_period[7] ));
 sky130_fd_sc_hd__dfrtp_2 _10882_ (.CLK(clknet_1_1__leaf__04675_),
    .D(net1429),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_clk_period[8] ));
 sky130_fd_sc_hd__dfrtp_2 _10883_ (.CLK(clknet_1_1__leaf__04675_),
    .D(net1423),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_clk_period[9] ));
 sky130_fd_sc_hd__dfrtp_2 _10884_ (.CLK(clknet_1_0__leaf__04675_),
    .D(net1291),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_th0_period[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10885_ (.CLK(clknet_1_1__leaf__04675_),
    .D(net1647),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_th0_period[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10886_ (.CLK(clknet_1_1__leaf__04675_),
    .D(net1640),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_th0_period[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10887_ (.CLK(clknet_1_0__leaf__04675_),
    .D(net1632),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th0_period[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10888_ (.CLK(clknet_1_0__leaf__04675_),
    .D(net1625),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th0_period[4] ));
 sky130_fd_sc_hd__dfrtp_2 _10889_ (.CLK(clknet_1_0__leaf__04675_),
    .D(net1618),
    .RESET_B(net1025),
    .Q(\u_ws281x.cfg_th0_period[5] ));
 sky130_fd_sc_hd__dfrtp_1 _10890_ (.CLK(clknet_1_1__leaf__04670_),
    .D(net1429),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_reset_period[8] ));
 sky130_fd_sc_hd__dfrtp_2 _10891_ (.CLK(clknet_1_1__leaf__04670_),
    .D(net1423),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_reset_period[9] ));
 sky130_fd_sc_hd__dfrtp_2 _10892_ (.CLK(clknet_1_0__leaf__04670_),
    .D(net1291),
    .RESET_B(net1022),
    .Q(\u_ws281x.cfg_reset_period[10] ));
 sky130_fd_sc_hd__dfrtp_1 _10893_ (.CLK(clknet_1_1__leaf__04670_),
    .D(net1647),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_reset_period[11] ));
 sky130_fd_sc_hd__dfrtp_1 _10894_ (.CLK(clknet_1_0__leaf__04670_),
    .D(net1640),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_reset_period[12] ));
 sky130_fd_sc_hd__dfrtp_1 _10895_ (.CLK(clknet_1_1__leaf__04670_),
    .D(net1632),
    .RESET_B(net1030),
    .Q(\u_ws281x.cfg_reset_period[13] ));
 sky130_fd_sc_hd__dfrtp_4 _10896_ (.CLK(clknet_1_0__leaf__04670_),
    .D(net1625),
    .RESET_B(net1023),
    .Q(\u_ws281x.cfg_reset_period[14] ));
 sky130_fd_sc_hd__dfrtp_1 _10897_ (.CLK(clknet_1_0__leaf__04670_),
    .D(net1618),
    .RESET_B(net1028),
    .Q(\u_ws281x.cfg_reset_period[15] ));
 sky130_fd_sc_hd__dfrtp_2 _10898_ (.CLK(clknet_1_0__leaf__04671_),
    .D(net1302),
    .RESET_B(net1031),
    .Q(\u_ws281x.cfg_reset_period[0] ));
 sky130_fd_sc_hd__dfrtp_1 _10899_ (.CLK(clknet_1_0__leaf__04671_),
    .D(net1576),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[1] ));
 sky130_fd_sc_hd__dfrtp_2 _10900_ (.CLK(clknet_1_0__leaf__04671_),
    .D(net1493),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[2] ));
 sky130_fd_sc_hd__dfrtp_2 _10901_ (.CLK(clknet_1_0__leaf__04671_),
    .D(net1470),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[3] ));
 sky130_fd_sc_hd__dfrtp_2 _10902_ (.CLK(clknet_1_1__leaf__04671_),
    .D(net1462),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[4] ));
 sky130_fd_sc_hd__dfrtp_1 _10903_ (.CLK(clknet_1_1__leaf__04671_),
    .D(net1453),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[5] ));
 sky130_fd_sc_hd__dfrtp_2 _10904_ (.CLK(clknet_1_1__leaf__04671_),
    .D(net1446),
    .RESET_B(net1034),
    .Q(\u_ws281x.cfg_reset_period[6] ));
 sky130_fd_sc_hd__dfrtp_1 _10905_ (.CLK(clknet_1_1__leaf__04671_),
    .D(net1437),
    .RESET_B(net1033),
    .Q(\u_ws281x.cfg_reset_period[7] ));
 sky130_fd_sc_hd__dfrtp_1 _10906_ (.CLK(_04666_),
    .D(net1302),
    .RESET_B(net1031),
    .Q(\u_ws281x.port0_enb ));
 sky130_fd_sc_hd__dfrtp_2 _10907_ (.CLK(_04667_),
    .D(net1576),
    .RESET_B(net1031),
    .Q(\u_ws281x.port1_enb ));
 sky130_fd_sc_hd__dfrtp_1 _10908_ (.CLK(_04668_),
    .D(net1493),
    .RESET_B(net1031),
    .Q(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10909_ (.CLK(_04669_),
    .D(net1470),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[3].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _10910_ (.CLK(_04660_),
    .D(_04345_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.wr_ptr ));
 sky130_fd_sc_hd__dfrtp_1 _10911_ (.CLK(_04661_),
    .D(_04346_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.rd_ptr ));
 sky130_fd_sc_hd__dfstp_2 _10912_ (.CLK(_04662_),
    .D(_00587_),
    .SET_B(net1036),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ));
 sky130_fd_sc_hd__dfrtp_2 _10913_ (.CLK(_04663_),
    .D(_00588_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.full ));
 sky130_fd_sc_hd__dfxtp_1 _10914_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1302),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10915_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1576),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10916_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1493),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10917_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1470),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10918_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1462),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10919_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1453),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10920_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1446),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10921_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1437),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10922_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1429),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10923_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1423),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10924_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1291),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10925_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1647),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10926_ (.CLK(clknet_1_1__leaf__04664_),
    .D(net1640),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10927_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1632),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10928_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1625),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10929_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1618),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10930_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1609),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10931_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1601),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10932_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1591),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10933_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1583),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10934_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1570),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10935_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1563),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10936_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1554),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10937_ (.CLK(clknet_1_0__leaf__04664_),
    .D(net1546),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10938_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1303),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10939_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1578),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10940_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1493),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10941_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1470),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10942_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1462),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10943_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1453),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10944_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1446),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10945_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1437),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10946_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1429),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10947_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1423),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10948_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1291),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10949_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1647),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10950_ (.CLK(clknet_1_1__leaf__04665_),
    .D(net1640),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10951_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1632),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10952_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1625),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10953_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1620),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10954_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1609),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10955_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1601),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10956_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1591),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10957_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1585),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10958_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1570),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10959_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1563),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10960_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1554),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10961_ (.CLK(clknet_1_0__leaf__04665_),
    .D(net1548),
    .Q(\u_ws281x.u_reg.gfifo[1].u_fifo.mem[0][23] ));
 sky130_fd_sc_hd__dfrtp_1 _10962_ (.CLK(_04654_),
    .D(_04343_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.wr_ptr ));
 sky130_fd_sc_hd__dfrtp_1 _10963_ (.CLK(_04655_),
    .D(_04344_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.rd_ptr ));
 sky130_fd_sc_hd__dfstp_2 _10964_ (.CLK(_04656_),
    .D(_00580_),
    .SET_B(net1021),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.empty ));
 sky130_fd_sc_hd__dfrtp_1 _10965_ (.CLK(_04657_),
    .D(_00581_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.full ));
 sky130_fd_sc_hd__dfxtp_1 _10966_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1303),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10967_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1578),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10968_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1493),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10969_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1472),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10970_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1464),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10971_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1453),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10972_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1447),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10973_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1439),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10974_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1429),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10975_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1423),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][9] ));
 sky130_fd_sc_hd__dfxtp_1 _10976_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1291),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][10] ));
 sky130_fd_sc_hd__dfxtp_1 _10977_ (.CLK(clknet_1_1__leaf__04658_),
    .D(net1647),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][11] ));
 sky130_fd_sc_hd__dfxtp_1 _10978_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1640),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][12] ));
 sky130_fd_sc_hd__dfxtp_1 _10979_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1632),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][13] ));
 sky130_fd_sc_hd__dfxtp_1 _10980_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1625),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][14] ));
 sky130_fd_sc_hd__dfxtp_1 _10981_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1620),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][15] ));
 sky130_fd_sc_hd__dfxtp_1 _10982_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1609),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][16] ));
 sky130_fd_sc_hd__dfxtp_1 _10983_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1601),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][17] ));
 sky130_fd_sc_hd__dfxtp_1 _10984_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1593),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][18] ));
 sky130_fd_sc_hd__dfxtp_1 _10985_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1583),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][19] ));
 sky130_fd_sc_hd__dfxtp_1 _10986_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1568),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][20] ));
 sky130_fd_sc_hd__dfxtp_1 _10987_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1561),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][21] ));
 sky130_fd_sc_hd__dfxtp_1 _10988_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1553),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][22] ));
 sky130_fd_sc_hd__dfxtp_1 _10989_ (.CLK(clknet_1_0__leaf__04658_),
    .D(net1548),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[1][23] ));
 sky130_fd_sc_hd__dfxtp_1 _10990_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1303),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][0] ));
 sky130_fd_sc_hd__dfxtp_1 _10991_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1578),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][1] ));
 sky130_fd_sc_hd__dfxtp_1 _10992_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1495),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][2] ));
 sky130_fd_sc_hd__dfxtp_1 _10993_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1472),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][3] ));
 sky130_fd_sc_hd__dfxtp_1 _10994_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1464),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][4] ));
 sky130_fd_sc_hd__dfxtp_1 _10995_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1455),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][5] ));
 sky130_fd_sc_hd__dfxtp_1 _10996_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1447),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][6] ));
 sky130_fd_sc_hd__dfxtp_1 _10997_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1439),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][7] ));
 sky130_fd_sc_hd__dfxtp_1 _10998_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1429),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][8] ));
 sky130_fd_sc_hd__dfxtp_1 _10999_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1423),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][9] ));
 sky130_fd_sc_hd__dfxtp_1 _11000_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1291),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][10] ));
 sky130_fd_sc_hd__dfxtp_1 _11001_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1647),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][11] ));
 sky130_fd_sc_hd__dfxtp_1 _11002_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1640),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][12] ));
 sky130_fd_sc_hd__dfxtp_1 _11003_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1632),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][13] ));
 sky130_fd_sc_hd__dfxtp_1 _11004_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1625),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][14] ));
 sky130_fd_sc_hd__dfxtp_1 _11005_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1620),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][15] ));
 sky130_fd_sc_hd__dfxtp_1 _11006_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1609),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][16] ));
 sky130_fd_sc_hd__dfxtp_1 _11007_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1601),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][17] ));
 sky130_fd_sc_hd__dfxtp_1 _11008_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1593),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][18] ));
 sky130_fd_sc_hd__dfxtp_1 _11009_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1583),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][19] ));
 sky130_fd_sc_hd__dfxtp_1 _11010_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1568),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][20] ));
 sky130_fd_sc_hd__dfxtp_1 _11011_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1561),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][21] ));
 sky130_fd_sc_hd__dfxtp_1 _11012_ (.CLK(clknet_1_0__leaf__04659_),
    .D(net1553),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][22] ));
 sky130_fd_sc_hd__dfxtp_1 _11013_ (.CLK(clknet_1_1__leaf__04659_),
    .D(net1548),
    .Q(\u_ws281x.u_reg.gfifo[0].u_fifo.mem[0][23] ));
 sky130_fd_sc_hd__dfrtp_4 _11014_ (.CLK(clknet_leaf_70_mclk),
    .D(_04681_),
    .RESET_B(net1032),
    .Q(\u_ws281x.u_txd_0.state ));
 sky130_fd_sc_hd__dfrtp_1 _11015_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00622_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11016_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00633_),
    .RESET_B(net1023),
    .Q(\u_ws281x.u_txd_0.led_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11017_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00638_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11018_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00639_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11019_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00640_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11020_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00641_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11021_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00642_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11022_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00643_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_txd_0.led_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11023_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00644_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_txd_0.led_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11024_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00645_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_txd_0.led_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11025_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00623_),
    .RESET_B(net1021),
    .Q(\u_ws281x.u_txd_0.led_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11026_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00624_),
    .RESET_B(net1022),
    .Q(\u_ws281x.u_txd_0.led_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11027_ (.CLK(clknet_1_1__leaf__04680_),
    .D(_00625_),
    .RESET_B(net1020),
    .Q(\u_ws281x.u_txd_0.led_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11028_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00626_),
    .RESET_B(net1020),
    .Q(\u_ws281x.u_txd_0.led_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11029_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00627_),
    .RESET_B(net1020),
    .Q(\u_ws281x.u_txd_0.led_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11030_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00628_),
    .RESET_B(net1020),
    .Q(\u_ws281x.u_txd_0.led_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11031_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00629_),
    .RESET_B(net1020),
    .Q(\u_ws281x.u_txd_0.led_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11032_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00630_),
    .RESET_B(net1019),
    .Q(\u_ws281x.u_txd_0.led_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11033_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00631_),
    .RESET_B(net1018),
    .Q(\u_ws281x.u_txd_0.led_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11034_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00632_),
    .RESET_B(net1018),
    .Q(\u_ws281x.u_txd_0.led_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11035_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00634_),
    .RESET_B(net1023),
    .Q(\u_ws281x.u_txd_0.led_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11036_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00635_),
    .RESET_B(net1018),
    .Q(\u_ws281x.u_txd_0.led_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11037_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00636_),
    .RESET_B(net1018),
    .Q(\u_ws281x.u_txd_0.led_data[22] ));
 sky130_fd_sc_hd__dfrtp_2 _11038_ (.CLK(clknet_1_0__leaf__04680_),
    .D(_00637_),
    .RESET_B(net1018),
    .Q(\u_ws281x.u_txd_0.led_data[23] ));
 sky130_fd_sc_hd__dfrtp_2 _11039_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00605_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_0.clk_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11040_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00612_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_0.clk_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11041_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00613_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_0.clk_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11042_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00614_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11043_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00615_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11044_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00616_),
    .RESET_B(net1035),
    .Q(\u_ws281x.u_txd_0.clk_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11045_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00617_),
    .RESET_B(net1035),
    .Q(\u_ws281x.u_txd_0.clk_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11046_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00618_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_0.clk_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11047_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00619_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_0.clk_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11048_ (.CLK(clknet_1_1__leaf__04679_),
    .D(_00620_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_0.clk_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11049_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00606_),
    .RESET_B(net1035),
    .Q(\u_ws281x.u_txd_0.clk_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11050_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00607_),
    .RESET_B(net1035),
    .Q(\u_ws281x.u_txd_0.clk_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11051_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00608_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11052_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00609_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11053_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00610_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11054_ (.CLK(clknet_1_0__leaf__04679_),
    .D(_00611_),
    .RESET_B(net1034),
    .Q(\u_ws281x.u_txd_0.clk_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11055_ (.CLK(_04678_),
    .D(_00621_),
    .RESET_B(net1031),
    .Q(\u_ws281x.port0_rd ));
 sky130_fd_sc_hd__dfrtp_1 _11056_ (.CLK(_04677_),
    .D(_00646_),
    .RESET_B(net1032),
    .Q(\u_ws281x.u_txd_0.txd ));
 sky130_fd_sc_hd__dfstp_1 _11057_ (.CLK(clknet_1_1__leaf__04676_),
    .D(_00600_),
    .SET_B(net1035),
    .Q(\u_ws281x.u_txd_0.bit_cnt[0] ));
 sky130_fd_sc_hd__dfstp_1 _11058_ (.CLK(clknet_1_1__leaf__04676_),
    .D(_00601_),
    .SET_B(net1035),
    .Q(\u_ws281x.u_txd_0.bit_cnt[1] ));
 sky130_fd_sc_hd__dfstp_1 _11059_ (.CLK(clknet_1_1__leaf__04676_),
    .D(_00602_),
    .SET_B(net1035),
    .Q(\u_ws281x.u_txd_0.bit_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11060_ (.CLK(clknet_1_0__leaf__04676_),
    .D(net2343),
    .RESET_B(net1032),
    .Q(\u_ws281x.u_txd_0.bit_cnt[3] ));
 sky130_fd_sc_hd__dfstp_1 _11061_ (.CLK(clknet_1_0__leaf__04676_),
    .D(_00604_),
    .SET_B(net1031),
    .Q(\u_ws281x.u_txd_0.bit_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11062_ (.CLK(clknet_leaf_69_mclk),
    .D(_04687_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.state ));
 sky130_fd_sc_hd__dfrtp_1 _11063_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00673_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.led_data[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11064_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00684_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.led_data[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11065_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00689_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11066_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00690_),
    .RESET_B(net1030),
    .Q(\u_ws281x.u_txd_1.led_data[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11067_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00691_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11068_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00692_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11069_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00693_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11070_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00694_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11071_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00695_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11072_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00696_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11073_ (.CLK(clknet_1_1__leaf__04686_),
    .D(_00674_),
    .RESET_B(net1029),
    .Q(\u_ws281x.u_txd_1.led_data[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11074_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00675_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11075_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00676_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11076_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00677_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11077_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00678_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11078_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00679_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11079_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00680_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11080_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00681_),
    .RESET_B(net1026),
    .Q(\u_ws281x.u_txd_1.led_data[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11081_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00682_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11082_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00683_),
    .RESET_B(net1026),
    .Q(\u_ws281x.u_txd_1.led_data[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11083_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00685_),
    .RESET_B(net1026),
    .Q(\u_ws281x.u_txd_1.led_data[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11084_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00686_),
    .RESET_B(net1026),
    .Q(\u_ws281x.u_txd_1.led_data[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11085_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00687_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11086_ (.CLK(clknet_1_0__leaf__04686_),
    .D(_00688_),
    .RESET_B(net1027),
    .Q(\u_ws281x.u_txd_1.led_data[23] ));
 sky130_fd_sc_hd__dfrtp_2 _11087_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00656_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_1.clk_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11088_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00663_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_1.clk_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11089_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00664_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_1.clk_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11090_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00665_),
    .RESET_B(net1037),
    .Q(\u_ws281x.u_txd_1.clk_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11091_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00666_),
    .RESET_B(net1037),
    .Q(\u_ws281x.u_txd_1.clk_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11092_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00667_),
    .RESET_B(net1037),
    .Q(\u_ws281x.u_txd_1.clk_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11093_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00668_),
    .RESET_B(net1037),
    .Q(\u_ws281x.u_txd_1.clk_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11094_ (.CLK(clknet_1_0__leaf__04685_),
    .D(_00669_),
    .RESET_B(net1037),
    .Q(\u_ws281x.u_txd_1.clk_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11095_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00670_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.clk_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11096_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00671_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11097_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00657_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11098_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00658_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11099_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00659_),
    .RESET_B(net1038),
    .Q(\u_ws281x.u_txd_1.clk_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11100_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00660_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11101_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00661_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11102_ (.CLK(clknet_1_1__leaf__04685_),
    .D(_00662_),
    .RESET_B(net1039),
    .Q(\u_ws281x.u_txd_1.clk_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11103_ (.CLK(_04684_),
    .D(_00672_),
    .RESET_B(net1036),
    .Q(\u_ws281x.port1_rd ));
 sky130_fd_sc_hd__dfrtp_1 _11104_ (.CLK(_04683_),
    .D(_00697_),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.txd ));
 sky130_fd_sc_hd__dfstp_1 _11105_ (.CLK(clknet_1_0__leaf__04682_),
    .D(_00651_),
    .SET_B(net1036),
    .Q(\u_ws281x.u_txd_1.bit_cnt[0] ));
 sky130_fd_sc_hd__dfstp_1 _11106_ (.CLK(clknet_1_1__leaf__04682_),
    .D(_00652_),
    .SET_B(net1037),
    .Q(\u_ws281x.u_txd_1.bit_cnt[1] ));
 sky130_fd_sc_hd__dfstp_1 _11107_ (.CLK(clknet_1_1__leaf__04682_),
    .D(_00653_),
    .SET_B(net1037),
    .Q(\u_ws281x.u_txd_1.bit_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11108_ (.CLK(clknet_1_0__leaf__04682_),
    .D(net2248),
    .RESET_B(net1036),
    .Q(\u_ws281x.u_txd_1.bit_cnt[3] ));
 sky130_fd_sc_hd__dfstp_1 _11109_ (.CLK(clknet_1_1__leaf__04682_),
    .D(_00655_),
    .SET_B(net1037),
    .Q(\u_ws281x.u_txd_1.bit_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11110_ (.CLK(clknet_1_1__leaf__04631_),
    .D(_00479_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11111_ (.CLK(clknet_1_0__leaf__04631_),
    .D(_00480_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11112_ (.CLK(clknet_1_0__leaf__04631_),
    .D(_00481_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11113_ (.CLK(clknet_1_1__leaf__04631_),
    .D(_00482_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11114_ (.CLK(clknet_1_1__leaf__04631_),
    .D(_00483_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11115_ (.CLK(clknet_1_1__leaf__04631_),
    .D(_00484_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11116_ (.CLK(clknet_1_1__leaf__04631_),
    .D(_00485_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11117_ (.CLK(clknet_1_0__leaf__04631_),
    .D(_00486_),
    .RESET_B(net967),
    .Q(\u_timer.u_pulse_1ms.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11118_ (.CLK(clknet_1_0__leaf__04631_),
    .D(_00487_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11119_ (.CLK(clknet_1_0__leaf__04631_),
    .D(_00488_),
    .RESET_B(net968),
    .Q(\u_timer.u_pulse_1ms.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11120_ (.CLK(clknet_1_1__leaf__04632_),
    .D(_00489_),
    .RESET_B(net759),
    .Q(\u_timer.u_pulse_1s.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11121_ (.CLK(clknet_1_1__leaf__04632_),
    .D(_00490_),
    .RESET_B(net759),
    .Q(\u_timer.u_pulse_1s.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11122_ (.CLK(clknet_1_1__leaf__04632_),
    .D(_00491_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11123_ (.CLK(clknet_1_0__leaf__04632_),
    .D(_00492_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11124_ (.CLK(clknet_1_0__leaf__04632_),
    .D(_00493_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11125_ (.CLK(clknet_1_0__leaf__04632_),
    .D(_00494_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11126_ (.CLK(clknet_1_0__leaf__04632_),
    .D(_00495_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11127_ (.CLK(clknet_1_0__leaf__04632_),
    .D(_00496_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11128_ (.CLK(clknet_1_1__leaf__04632_),
    .D(_00497_),
    .RESET_B(net759),
    .Q(\u_timer.u_pulse_1s.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11129_ (.CLK(clknet_1_1__leaf__04632_),
    .D(_00498_),
    .RESET_B(net758),
    .Q(\u_timer.u_pulse_1s.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11130_ (.CLK(clknet_leaf_47_mclk),
    .D(_00500_),
    .RESET_B(net969),
    .Q(\u_timer.u_pulse_1us.cnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11131_ (.CLK(clknet_leaf_47_mclk),
    .D(_00501_),
    .RESET_B(net969),
    .Q(\u_timer.u_pulse_1us.cnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11132_ (.CLK(clknet_leaf_47_mclk),
    .D(_00502_),
    .RESET_B(net974),
    .Q(\u_timer.u_pulse_1us.cnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11133_ (.CLK(clknet_leaf_48_mclk),
    .D(_00503_),
    .RESET_B(net974),
    .Q(\u_timer.u_pulse_1us.cnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11134_ (.CLK(clknet_leaf_48_mclk),
    .D(_00504_),
    .RESET_B(net974),
    .Q(\u_timer.u_pulse_1us.cnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11135_ (.CLK(clknet_leaf_48_mclk),
    .D(_00505_),
    .RESET_B(net974),
    .Q(\u_timer.u_pulse_1us.cnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11136_ (.CLK(clknet_leaf_48_mclk),
    .D(_00506_),
    .RESET_B(net974),
    .Q(\u_timer.u_pulse_1us.cnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11137_ (.CLK(clknet_leaf_48_mclk),
    .D(_00507_),
    .RESET_B(net973),
    .Q(\u_timer.u_pulse_1us.cnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11138_ (.CLK(clknet_leaf_48_mclk),
    .D(_00508_),
    .RESET_B(net973),
    .Q(\u_timer.u_pulse_1us.cnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11139_ (.CLK(clknet_leaf_48_mclk),
    .D(_00509_),
    .RESET_B(net973),
    .Q(\u_timer.u_pulse_1us.cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11140_ (.CLK(clknet_leaf_48_mclk),
    .D(_00499_),
    .RESET_B(net969),
    .Q(\u_gpio.pulse_1us ));
 sky130_fd_sc_hd__dfrtp_4 _11141_ (.CLK(clknet_leaf_55_mclk),
    .D(_00510_),
    .RESET_B(net930),
    .Q(\u_timer.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _11142_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[0] ),
    .RESET_B(net933),
    .Q(\u_timer.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11143_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[1] ),
    .RESET_B(net933),
    .Q(\u_timer.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11144_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[2] ),
    .RESET_B(net922),
    .Q(\u_timer.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11145_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[3] ),
    .RESET_B(net923),
    .Q(\u_timer.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11146_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[4] ),
    .RESET_B(net931),
    .Q(\u_timer.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11147_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[5] ),
    .RESET_B(net930),
    .Q(\u_timer.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11148_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[6] ),
    .RESET_B(net963),
    .Q(\u_timer.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11149_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[7] ),
    .RESET_B(net963),
    .Q(\u_timer.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11150_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[8] ),
    .RESET_B(net962),
    .Q(\u_timer.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11151_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[9] ),
    .RESET_B(net962),
    .Q(\u_timer.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11152_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[10] ),
    .RESET_B(net961),
    .Q(\u_timer.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11153_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[11] ),
    .RESET_B(net960),
    .Q(\u_timer.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11154_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[12] ),
    .RESET_B(net960),
    .Q(\u_timer.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11155_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[13] ),
    .RESET_B(net960),
    .Q(\u_timer.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11156_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[14] ),
    .RESET_B(net960),
    .Q(\u_timer.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11157_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[15] ),
    .RESET_B(net960),
    .Q(\u_timer.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11158_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[16] ),
    .RESET_B(net934),
    .Q(\u_timer.reg_rdata[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11159_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[17] ),
    .RESET_B(net934),
    .Q(\u_timer.reg_rdata[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11160_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[18] ),
    .RESET_B(net935),
    .Q(\u_timer.reg_rdata[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11161_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[19] ),
    .RESET_B(net931),
    .Q(\u_timer.reg_rdata[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11162_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[20] ),
    .RESET_B(net930),
    .Q(\u_timer.reg_rdata[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11163_ (.CLK(clknet_2_2__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[21] ),
    .RESET_B(net935),
    .Q(\u_timer.reg_rdata[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11164_ (.CLK(clknet_2_3__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[22] ),
    .RESET_B(net931),
    .Q(\u_timer.reg_rdata[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11165_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[23] ),
    .RESET_B(net931),
    .Q(\u_timer.reg_rdata[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11166_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[24] ),
    .RESET_B(net813),
    .Q(\u_timer.reg_rdata[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11167_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[25] ),
    .RESET_B(net810),
    .Q(\u_timer.reg_rdata[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11168_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[26] ),
    .RESET_B(net812),
    .Q(\u_timer.reg_rdata[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11169_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[27] ),
    .RESET_B(net921),
    .Q(\u_timer.reg_rdata[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11170_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[28] ),
    .RESET_B(net921),
    .Q(\u_timer.reg_rdata[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11171_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[29] ),
    .RESET_B(net810),
    .Q(\u_timer.reg_rdata[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11172_ (.CLK(clknet_2_0__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[30] ),
    .RESET_B(net809),
    .Q(\u_timer.reg_rdata[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11173_ (.CLK(clknet_2_1__leaf__04633_),
    .D(\u_timer.u_reg.reg_out[31] ),
    .RESET_B(net809),
    .Q(\u_timer.reg_rdata[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11174_ (.CLK(clknet_1_1__leaf__04646_),
    .D(net1606),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11175_ (.CLK(clknet_1_1__leaf__04646_),
    .D(net1599),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11176_ (.CLK(clknet_1_1__leaf__04646_),
    .D(net1590),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11177_ (.CLK(clknet_1_0__leaf__04646_),
    .D(net1581),
    .RESET_B(net925),
    .Q(\u_timer.u_reg.reg_3[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11178_ (.CLK(clknet_1_0__leaf__04646_),
    .D(net1568),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_3[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11179_ (.CLK(clknet_1_1__leaf__04646_),
    .D(net1561),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_3[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11180_ (.CLK(clknet_1_0__leaf__04646_),
    .D(net1553),
    .RESET_B(net925),
    .Q(\u_timer.u_reg.reg_3[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11181_ (.CLK(clknet_1_0__leaf__04646_),
    .D(net1546),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_3[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11182_ (.CLK(clknet_1_1__leaf__04647_),
    .D(net1538),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_3[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11183_ (.CLK(clknet_1_0__leaf__04647_),
    .D(net1530),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_3[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11184_ (.CLK(clknet_1_1__leaf__04647_),
    .D(net1524),
    .RESET_B(net922),
    .Q(\u_timer.u_reg.reg_3[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11185_ (.CLK(clknet_1_1__leaf__04647_),
    .D(net1517),
    .RESET_B(net922),
    .Q(\u_timer.u_reg.reg_3[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11186_ (.CLK(clknet_1_1__leaf__04647_),
    .D(net1508),
    .RESET_B(net921),
    .Q(\u_timer.u_reg.reg_3[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11187_ (.CLK(clknet_1_0__leaf__04647_),
    .D(net1500),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_3[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11188_ (.CLK(clknet_1_0__leaf__04647_),
    .D(net1484),
    .RESET_B(net808),
    .Q(\u_timer.u_reg.reg_3[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11189_ (.CLK(clknet_1_0__leaf__04647_),
    .D(net1478),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_3[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11190_ (.CLK(clknet_1_1__leaf__04648_),
    .D(net1302),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11191_ (.CLK(clknet_1_1__leaf__04648_),
    .D(net1576),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11192_ (.CLK(clknet_1_1__leaf__04648_),
    .D(net1495),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11193_ (.CLK(clknet_1_1__leaf__04648_),
    .D(net1472),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11194_ (.CLK(clknet_1_0__leaf__04648_),
    .D(net1462),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11195_ (.CLK(clknet_1_0__leaf__04648_),
    .D(net1454),
    .RESET_B(net959),
    .Q(\u_timer.cfg_timer2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11196_ (.CLK(clknet_1_0__leaf__04648_),
    .D(net1446),
    .RESET_B(net959),
    .Q(\u_timer.cfg_timer2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11197_ (.CLK(clknet_1_0__leaf__04648_),
    .D(net1437),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11198_ (.CLK(clknet_1_1__leaf__04649_),
    .D(net1429),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11199_ (.CLK(clknet_1_1__leaf__04649_),
    .D(net1423),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11200_ (.CLK(clknet_1_1__leaf__04649_),
    .D(net1291),
    .RESET_B(net956),
    .Q(\u_timer.cfg_timer2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11201_ (.CLK(clknet_1_1__leaf__04649_),
    .D(net1647),
    .RESET_B(net956),
    .Q(\u_timer.cfg_timer2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11202_ (.CLK(clknet_1_0__leaf__04649_),
    .D(net1640),
    .RESET_B(net956),
    .Q(\u_timer.cfg_timer2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11203_ (.CLK(clknet_1_0__leaf__04649_),
    .D(net1632),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11204_ (.CLK(clknet_1_0__leaf__04649_),
    .D(net1625),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11205_ (.CLK(clknet_1_0__leaf__04649_),
    .D(net1618),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11206_ (.CLK(clknet_1_1__leaf__04642_),
    .D(net1611),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11207_ (.CLK(clknet_1_1__leaf__04642_),
    .D(net1599),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11208_ (.CLK(clknet_1_1__leaf__04642_),
    .D(net1591),
    .RESET_B(net928),
    .Q(\u_timer.cfg_timer1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11209_ (.CLK(clknet_1_0__leaf__04642_),
    .D(net1582),
    .RESET_B(net929),
    .Q(\u_timer.u_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11210_ (.CLK(clknet_1_0__leaf__04642_),
    .D(net1568),
    .RESET_B(net932),
    .Q(\u_timer.u_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11211_ (.CLK(clknet_1_1__leaf__04642_),
    .D(net1561),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11212_ (.CLK(clknet_1_0__leaf__04642_),
    .D(net1553),
    .RESET_B(net928),
    .Q(\u_timer.u_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11213_ (.CLK(clknet_1_0__leaf__04642_),
    .D(net1546),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11214_ (.CLK(clknet_1_0__leaf__04643_),
    .D(net1538),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11215_ (.CLK(clknet_1_0__leaf__04643_),
    .D(net1530),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11216_ (.CLK(clknet_1_1__leaf__04643_),
    .D(net1523),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11217_ (.CLK(clknet_1_1__leaf__04643_),
    .D(net1516),
    .RESET_B(net921),
    .Q(\u_timer.u_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11218_ (.CLK(clknet_1_1__leaf__04643_),
    .D(net1509),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11219_ (.CLK(clknet_1_0__leaf__04643_),
    .D(net1500),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11220_ (.CLK(clknet_1_0__leaf__04643_),
    .D(net1484),
    .RESET_B(net808),
    .Q(\u_timer.u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11221_ (.CLK(clknet_1_1__leaf__04643_),
    .D(net1478),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11222_ (.CLK(clknet_1_1__leaf__04644_),
    .D(net1302),
    .RESET_B(net966),
    .Q(\u_timer.cfg_timer1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11223_ (.CLK(clknet_1_1__leaf__04644_),
    .D(net1576),
    .RESET_B(net966),
    .Q(\u_timer.cfg_timer1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11224_ (.CLK(clknet_1_1__leaf__04644_),
    .D(net1495),
    .RESET_B(net966),
    .Q(\u_timer.cfg_timer1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11225_ (.CLK(clknet_1_1__leaf__04644_),
    .D(net1472),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11226_ (.CLK(clknet_1_0__leaf__04644_),
    .D(net1462),
    .RESET_B(net965),
    .Q(\u_timer.cfg_timer1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11227_ (.CLK(clknet_1_0__leaf__04644_),
    .D(net1454),
    .RESET_B(net959),
    .Q(\u_timer.cfg_timer1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11228_ (.CLK(clknet_1_0__leaf__04644_),
    .D(net1446),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11229_ (.CLK(clknet_1_0__leaf__04644_),
    .D(net1437),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11230_ (.CLK(clknet_1_1__leaf__04645_),
    .D(net1429),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11231_ (.CLK(clknet_1_1__leaf__04645_),
    .D(net1423),
    .RESET_B(net958),
    .Q(\u_timer.cfg_timer1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11232_ (.CLK(clknet_1_1__leaf__04645_),
    .D(net1291),
    .RESET_B(net956),
    .Q(\u_timer.cfg_timer1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11233_ (.CLK(clknet_1_1__leaf__04645_),
    .D(net1647),
    .RESET_B(net956),
    .Q(\u_timer.cfg_timer1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11234_ (.CLK(clknet_1_0__leaf__04645_),
    .D(net1640),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11235_ (.CLK(clknet_1_0__leaf__04645_),
    .D(net1632),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11236_ (.CLK(clknet_1_0__leaf__04645_),
    .D(net1625),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11237_ (.CLK(clknet_1_0__leaf__04645_),
    .D(net1618),
    .RESET_B(net955),
    .Q(\u_timer.cfg_timer1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11238_ (.CLK(clknet_1_1__leaf__04638_),
    .D(net1607),
    .RESET_B(net934),
    .Q(\u_timer.cfg_timer0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11239_ (.CLK(clknet_1_1__leaf__04638_),
    .D(net1600),
    .RESET_B(net934),
    .Q(\u_timer.cfg_timer0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11240_ (.CLK(clknet_1_1__leaf__04638_),
    .D(net1591),
    .RESET_B(net933),
    .Q(\u_timer.cfg_timer0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11241_ (.CLK(clknet_1_0__leaf__04638_),
    .D(net1583),
    .RESET_B(net932),
    .Q(\u_timer.u_reg.reg_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11242_ (.CLK(clknet_1_0__leaf__04638_),
    .D(net1568),
    .RESET_B(net932),
    .Q(\u_timer.u_reg.reg_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11243_ (.CLK(clknet_1_1__leaf__04638_),
    .D(net1561),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11244_ (.CLK(clknet_1_0__leaf__04638_),
    .D(net1553),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11245_ (.CLK(clknet_1_0__leaf__04638_),
    .D(net1546),
    .RESET_B(net932),
    .Q(\u_timer.u_reg.reg_1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11246_ (.CLK(clknet_1_1__leaf__04639_),
    .D(net1538),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11247_ (.CLK(clknet_1_0__leaf__04639_),
    .D(net1530),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11248_ (.CLK(clknet_1_1__leaf__04639_),
    .D(net1524),
    .RESET_B(net921),
    .Q(\u_timer.u_reg.reg_1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11249_ (.CLK(clknet_1_1__leaf__04639_),
    .D(net1517),
    .RESET_B(net922),
    .Q(\u_timer.u_reg.reg_1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11250_ (.CLK(clknet_1_1__leaf__04639_),
    .D(net1509),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11251_ (.CLK(clknet_1_0__leaf__04639_),
    .D(net1500),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11252_ (.CLK(clknet_1_0__leaf__04639_),
    .D(net1484),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11253_ (.CLK(clknet_1_0__leaf__04639_),
    .D(net1478),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11254_ (.CLK(clknet_1_1__leaf__04640_),
    .D(net1302),
    .RESET_B(net970),
    .Q(\u_timer.cfg_timer0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11255_ (.CLK(clknet_1_1__leaf__04640_),
    .D(net1576),
    .RESET_B(net970),
    .Q(\u_timer.cfg_timer0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11256_ (.CLK(clknet_1_1__leaf__04640_),
    .D(net1495),
    .RESET_B(net970),
    .Q(\u_timer.cfg_timer0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11257_ (.CLK(clknet_1_1__leaf__04640_),
    .D(net1472),
    .RESET_B(net971),
    .Q(\u_timer.cfg_timer0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11258_ (.CLK(clknet_1_0__leaf__04640_),
    .D(net1462),
    .RESET_B(net970),
    .Q(\u_timer.cfg_timer0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11259_ (.CLK(clknet_1_0__leaf__04640_),
    .D(net1455),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11260_ (.CLK(clknet_1_0__leaf__04640_),
    .D(net1446),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11261_ (.CLK(clknet_1_0__leaf__04640_),
    .D(net1437),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11262_ (.CLK(clknet_1_1__leaf__04641_),
    .D(net1431),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11263_ (.CLK(clknet_1_1__leaf__04641_),
    .D(net1424),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11264_ (.CLK(clknet_1_1__leaf__04641_),
    .D(net1292),
    .RESET_B(net963),
    .Q(\u_timer.cfg_timer0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11265_ (.CLK(clknet_1_1__leaf__04641_),
    .D(net1649),
    .RESET_B(net962),
    .Q(\u_timer.cfg_timer0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11266_ (.CLK(clknet_1_0__leaf__04641_),
    .D(net1640),
    .RESET_B(net961),
    .Q(\u_timer.cfg_timer0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11267_ (.CLK(clknet_1_0__leaf__04641_),
    .D(net1634),
    .RESET_B(net964),
    .Q(\u_timer.cfg_timer0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11268_ (.CLK(clknet_1_0__leaf__04641_),
    .D(net1625),
    .RESET_B(net961),
    .Q(\u_timer.cfg_timer0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11269_ (.CLK(clknet_1_0__leaf__04641_),
    .D(net1618),
    .RESET_B(net961),
    .Q(\u_timer.cfg_timer0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11270_ (.CLK(clknet_1_1__leaf__04634_),
    .D(net1607),
    .RESET_B(net934),
    .Q(\u_timer.u_reg.reg_0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11271_ (.CLK(clknet_1_1__leaf__04634_),
    .D(net1600),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11272_ (.CLK(clknet_1_1__leaf__04634_),
    .D(net1591),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11273_ (.CLK(clknet_1_0__leaf__04634_),
    .D(net1583),
    .RESET_B(net932),
    .Q(\u_timer.u_reg.reg_0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11274_ (.CLK(clknet_1_0__leaf__04634_),
    .D(net1568),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11275_ (.CLK(clknet_1_1__leaf__04634_),
    .D(net1561),
    .RESET_B(net933),
    .Q(\u_timer.u_reg.reg_0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11276_ (.CLK(clknet_1_0__leaf__04634_),
    .D(net1553),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11277_ (.CLK(clknet_1_0__leaf__04634_),
    .D(net1546),
    .RESET_B(net930),
    .Q(\u_timer.u_reg.reg_0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11278_ (.CLK(clknet_1_1__leaf__04635_),
    .D(net1538),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11279_ (.CLK(clknet_1_0__leaf__04635_),
    .D(net1530),
    .RESET_B(net812),
    .Q(\u_timer.u_reg.reg_0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11280_ (.CLK(clknet_1_1__leaf__04635_),
    .D(net1523),
    .RESET_B(net813),
    .Q(\u_timer.u_reg.reg_0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11281_ (.CLK(clknet_1_1__leaf__04635_),
    .D(net1516),
    .RESET_B(net921),
    .Q(\u_timer.u_reg.reg_0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11282_ (.CLK(clknet_1_1__leaf__04635_),
    .D(net1509),
    .RESET_B(net921),
    .Q(\u_timer.u_reg.reg_0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11283_ (.CLK(clknet_1_0__leaf__04635_),
    .D(net1501),
    .RESET_B(net810),
    .Q(\u_timer.u_reg.reg_0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11284_ (.CLK(clknet_1_0__leaf__04635_),
    .D(net1485),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11285_ (.CLK(clknet_1_0__leaf__04635_),
    .D(net1478),
    .RESET_B(net809),
    .Q(\u_timer.u_reg.reg_0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11286_ (.CLK(clknet_1_1__leaf__04636_),
    .D(net1302),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11287_ (.CLK(clknet_1_1__leaf__04636_),
    .D(net1576),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11288_ (.CLK(clknet_1_1__leaf__04636_),
    .D(net1495),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11289_ (.CLK(clknet_1_0__leaf__04636_),
    .D(net1472),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11290_ (.CLK(clknet_1_0__leaf__04636_),
    .D(net1462),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11291_ (.CLK(clknet_1_1__leaf__04636_),
    .D(net1454),
    .RESET_B(net970),
    .Q(\u_timer.cfg_pulse_1us[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11292_ (.CLK(clknet_1_0__leaf__04636_),
    .D(net1446),
    .RESET_B(net972),
    .Q(\u_timer.cfg_pulse_1us[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11293_ (.CLK(clknet_1_0__leaf__04636_),
    .D(net1437),
    .RESET_B(net972),
    .Q(\u_timer.cfg_pulse_1us[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11294_ (.CLK(clknet_1_1__leaf__04637_),
    .D(net1429),
    .RESET_B(net962),
    .Q(\u_timer.cfg_pulse_1us[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11295_ (.CLK(clknet_1_1__leaf__04637_),
    .D(net1423),
    .RESET_B(net962),
    .Q(\u_timer.cfg_pulse_1us[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11296_ (.CLK(clknet_1_1__leaf__04637_),
    .D(net1291),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11297_ (.CLK(clknet_1_1__leaf__04637_),
    .D(net1647),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11298_ (.CLK(clknet_1_0__leaf__04637_),
    .D(net1642),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11299_ (.CLK(clknet_1_0__leaf__04637_),
    .D(net1632),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11300_ (.CLK(clknet_1_0__leaf__04637_),
    .D(net1627),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11301_ (.CLK(clknet_1_0__leaf__04637_),
    .D(net1618),
    .RESET_B(net961),
    .Q(\u_timer.u_reg.reg_0[15] ));
 sky130_fd_sc_hd__dfstp_1 _11302_ (.CLK(clknet_leaf_54_mclk),
    .D(\u_timer.u_timer_0.timer_hit ),
    .SET_B(net934),
    .Q(\u_timer.u_timer_0.timer_hit_s1 ));
 sky130_fd_sc_hd__dfrtp_1 _11303_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00527_),
    .RESET_B(net971),
    .Q(\u_timer.u_timer_0.timer_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11304_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00534_),
    .RESET_B(net971),
    .Q(\u_timer.u_timer_0.timer_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11305_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00535_),
    .RESET_B(net971),
    .Q(\u_timer.u_timer_0.timer_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11306_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00536_),
    .RESET_B(net972),
    .Q(\u_timer.u_timer_0.timer_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11307_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00537_),
    .RESET_B(net971),
    .Q(\u_timer.u_timer_0.timer_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11308_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00538_),
    .RESET_B(net971),
    .Q(\u_timer.u_timer_0.timer_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11309_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00539_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11310_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00540_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11311_ (.CLK(clknet_1_1__leaf__04650_),
    .D(_00541_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11312_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00542_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11313_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00528_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11314_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00529_),
    .RESET_B(net963),
    .Q(\u_timer.u_timer_0.timer_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11315_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00530_),
    .RESET_B(net960),
    .Q(\u_timer.u_timer_0.timer_counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11316_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00531_),
    .RESET_B(net960),
    .Q(\u_timer.u_timer_0.timer_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11317_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00532_),
    .RESET_B(net960),
    .Q(\u_timer.u_timer_0.timer_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11318_ (.CLK(clknet_1_0__leaf__04650_),
    .D(_00533_),
    .RESET_B(net960),
    .Q(\u_timer.u_timer_0.timer_counter[15] ));
 sky130_fd_sc_hd__dfstp_1 _11319_ (.CLK(clknet_leaf_53_mclk),
    .D(\u_timer.u_timer_1.timer_hit ),
    .SET_B(net928),
    .Q(\u_timer.u_timer_1.timer_hit_s1 ));
 sky130_fd_sc_hd__dfrtp_1 _11320_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00544_),
    .RESET_B(net966),
    .Q(\u_timer.u_timer_1.timer_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11321_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00551_),
    .RESET_B(net966),
    .Q(\u_timer.u_timer_1.timer_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11322_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00552_),
    .RESET_B(net966),
    .Q(\u_timer.u_timer_1.timer_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11323_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00553_),
    .RESET_B(net965),
    .Q(\u_timer.u_timer_1.timer_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11324_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00554_),
    .RESET_B(net965),
    .Q(\u_timer.u_timer_1.timer_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11325_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00555_),
    .RESET_B(net965),
    .Q(\u_timer.u_timer_1.timer_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11326_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00556_),
    .RESET_B(net959),
    .Q(\u_timer.u_timer_1.timer_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11327_ (.CLK(clknet_1_1__leaf__04651_),
    .D(_00557_),
    .RESET_B(net958),
    .Q(\u_timer.u_timer_1.timer_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11328_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00558_),
    .RESET_B(net958),
    .Q(\u_timer.u_timer_1.timer_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11329_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00559_),
    .RESET_B(net958),
    .Q(\u_timer.u_timer_1.timer_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11330_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00545_),
    .RESET_B(net956),
    .Q(\u_timer.u_timer_1.timer_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11331_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00546_),
    .RESET_B(net956),
    .Q(\u_timer.u_timer_1.timer_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11332_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00547_),
    .RESET_B(net955),
    .Q(\u_timer.u_timer_1.timer_counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11333_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00548_),
    .RESET_B(net955),
    .Q(\u_timer.u_timer_1.timer_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11334_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00549_),
    .RESET_B(net955),
    .Q(\u_timer.u_timer_1.timer_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11335_ (.CLK(clknet_1_0__leaf__04651_),
    .D(_00550_),
    .RESET_B(net929),
    .Q(\u_timer.u_timer_1.timer_counter[15] ));
 sky130_fd_sc_hd__dfstp_1 _11336_ (.CLK(clknet_leaf_53_mclk),
    .D(\u_timer.u_timer_2.timer_hit ),
    .SET_B(net927),
    .Q(\u_timer.u_timer_2.timer_hit_s1 ));
 sky130_fd_sc_hd__dfrtp_1 _11337_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00561_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11338_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00568_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11339_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00569_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11340_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00570_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11341_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00571_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11342_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00572_),
    .RESET_B(net967),
    .Q(\u_timer.u_timer_2.timer_counter[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11343_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00573_),
    .RESET_B(net959),
    .Q(\u_timer.u_timer_2.timer_counter[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11344_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00574_),
    .RESET_B(net959),
    .Q(\u_timer.u_timer_2.timer_counter[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11345_ (.CLK(clknet_1_1__leaf__04652_),
    .D(_00575_),
    .RESET_B(net959),
    .Q(\u_timer.u_timer_2.timer_counter[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11346_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00576_),
    .RESET_B(net959),
    .Q(\u_timer.u_timer_2.timer_counter[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11347_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00562_),
    .RESET_B(net957),
    .Q(\u_timer.u_timer_2.timer_counter[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11348_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00563_),
    .RESET_B(net957),
    .Q(\u_timer.u_timer_2.timer_counter[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11349_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00564_),
    .RESET_B(net957),
    .Q(\u_timer.u_timer_2.timer_counter[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11350_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00565_),
    .RESET_B(net957),
    .Q(\u_timer.u_timer_2.timer_counter[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11351_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00566_),
    .RESET_B(net957),
    .Q(\u_timer.u_timer_2.timer_counter[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11352_ (.CLK(clknet_1_0__leaf__04652_),
    .D(_00567_),
    .RESET_B(net928),
    .Q(\u_timer.u_timer_2.timer_counter[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11353_ (.CLK(clknet_1_0__leaf__04629_),
    .D(_00762_),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11354_ (.CLK(clknet_1_0__leaf__04629_),
    .D(_00763_),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11355_ (.CLK(clknet_1_0__leaf__04629_),
    .D(_00764_),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11356_ (.CLK(clknet_1_0__leaf__04629_),
    .D(_00765_),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11357_ (.CLK(clknet_1_1__leaf__04629_),
    .D(_00766_),
    .RESET_B(net934),
    .Q(\u_semaphore.reg_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11358_ (.CLK(clknet_1_1__leaf__04629_),
    .D(_00767_),
    .RESET_B(net934),
    .Q(\u_semaphore.reg_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11359_ (.CLK(clknet_1_1__leaf__04629_),
    .D(_00768_),
    .RESET_B(net934),
    .Q(\u_semaphore.reg_0[14] ));
 sky130_fd_sc_hd__dfrtp_2 _11360_ (.CLK(clknet_1_1__leaf__04629_),
    .D(_00769_),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_0[15] ));
 sky130_fd_sc_hd__dfxtp_1 _11361_ (.CLK(clknet_1_1__leaf__04419_),
    .D(_00770_),
    .Q(\u_glbl_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfxtp_1 _11362_ (.CLK(clknet_1_1__leaf__04419_),
    .D(_00771_),
    .Q(\u_glbl_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfxtp_1 _11363_ (.CLK(clknet_1_0__leaf__04419_),
    .D(_00772_),
    .Q(\u_glbl_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfxtp_1 _11364_ (.CLK(clknet_1_0__leaf__04419_),
    .D(_00773_),
    .Q(\u_glbl_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfxtp_1 _11365_ (.CLK(clknet_1_0__leaf__04419_),
    .D(_00774_),
    .Q(\u_glbl_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfxtp_1 _11366_ (.CLK(clknet_1_0__leaf__04419_),
    .D(_00775_),
    .Q(\u_glbl_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11367_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[0] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11368_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[1] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11369_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[2] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11370_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[3] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11371_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[4] ),
    .RESET_B(net980),
    .Q(\u_semaphore.reg_rdata[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11372_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[5] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11373_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[6] ),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_rdata[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11374_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[7] ),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_rdata[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11375_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[8] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11376_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[9] ),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_rdata[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11377_ (.CLK(clknet_1_0__leaf__04628_),
    .D(\u_semaphore.reg_out[10] ),
    .RESET_B(net978),
    .Q(\u_semaphore.reg_rdata[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11378_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[11] ),
    .RESET_B(net1018),
    .Q(\u_semaphore.reg_rdata[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11379_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[12] ),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_rdata[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11380_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[13] ),
    .RESET_B(net992),
    .Q(\u_semaphore.reg_rdata[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11381_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[14] ),
    .RESET_B(net1018),
    .Q(\u_semaphore.reg_rdata[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11382_ (.CLK(clknet_1_1__leaf__04628_),
    .D(\u_semaphore.reg_out[15] ),
    .RESET_B(net960),
    .Q(\u_semaphore.reg_rdata[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11383_ (.CLK(clknet_leaf_55_mclk),
    .D(_00476_),
    .RESET_B(net931),
    .Q(\u_semaphore.reg_ack ));
 sky130_fd_sc_hd__dfrtp_1 _11384_ (.CLK(clknet_4_0__leaf_mclk),
    .D(net1690),
    .RESET_B(net134),
    .Q(\u_rst_sync.in_data_s ));
 sky130_fd_sc_hd__conb_1 _11384__1690 (.HI(net1690));
 sky130_fd_sc_hd__dfrtp_1 _11385_ (.CLK(clknet_leaf_118_mclk),
    .D(net2054),
    .RESET_B(net134),
    .Q(\u_rst_sync.in_data_2s ));
 sky130_fd_sc_hd__dfrtp_1 _11386_ (.CLK(clknet_leaf_76_mclk),
    .D(_00308_),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_run ));
 sky130_fd_sc_hd__dfrtp_1 _11387_ (.CLK(clknet_leaf_87_mclk),
    .D(_00309_),
    .RESET_B(net889),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_run ));
 sky130_fd_sc_hd__dfrtp_4 _11388_ (.CLK(clknet_leaf_96_mclk),
    .D(_00310_),
    .RESET_B(net844),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_run ));
 sky130_fd_sc_hd__dfrtp_2 _11389_ (.CLK(clknet_leaf_79_mclk),
    .D(_00311_),
    .RESET_B(net976),
    .Q(\u_pwm.reg_ack_glbl ));
 sky130_fd_sc_hd__dfrtp_1 _11390_ (.CLK(clknet_1_0__leaf__04552_),
    .D(net1605),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_dupdate ));
 sky130_fd_sc_hd__dfrtp_1 _11391_ (.CLK(clknet_1_1__leaf__04552_),
    .D(net1596),
    .RESET_B(net877),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_dupdate ));
 sky130_fd_sc_hd__dfrtp_1 _11392_ (.CLK(clknet_1_0__leaf__04552_),
    .D(net1588),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_dupdate ));
 sky130_fd_sc_hd__dfrtp_4 _11393_ (.CLK(clknet_1_1__leaf__04551_),
    .D(net1296),
    .RESET_B(net877),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_enb ));
 sky130_fd_sc_hd__dfrtp_4 _11394_ (.CLK(clknet_1_0__leaf__04551_),
    .D(net1574),
    .RESET_B(net877),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_enb ));
 sky130_fd_sc_hd__dfrtp_4 _11395_ (.CLK(clknet_1_0__leaf__04551_),
    .D(net1490),
    .RESET_B(net877),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_enb ));
 sky130_fd_sc_hd__dfrtp_1 _11396_ (.CLK(_04556_),
    .D(net1297),
    .RESET_B(net888),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11397_ (.CLK(_04557_),
    .D(net1574),
    .RESET_B(net889),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11398_ (.CLK(_04558_),
    .D(net1491),
    .RESET_B(net876),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11399_ (.CLK(_04559_),
    .D(net1470),
    .RESET_B(net1000),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[3].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11400_ (.CLK(_04560_),
    .D(net1461),
    .RESET_B(net1000),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[4].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11401_ (.CLK(_04561_),
    .D(net1453),
    .RESET_B(net1000),
    .Q(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[5].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11402_ (.CLK(_04553_),
    .D(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.hware_req ),
    .RESET_B(net999),
    .Q(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11403_ (.CLK(_04554_),
    .D(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.hware_req ),
    .RESET_B(net889),
    .Q(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[1].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11404_ (.CLK(_04555_),
    .D(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.hware_req ),
    .RESET_B(net876),
    .Q(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ));
 sky130_fd_sc_hd__dfrtp_1 _11405_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2174),
    .RESET_B(net1009),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_scale[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11406_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2157),
    .RESET_B(net1009),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_scale[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11407_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2184),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_scale[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11408_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2165),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_scale[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11409_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2166),
    .RESET_B(net1001),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_oneshot ));
 sky130_fd_sc_hd__dfrtp_1 _11410_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2193),
    .RESET_B(net1000),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_gpio_enb ));
 sky130_fd_sc_hd__dfrtp_1 _11411_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2187),
    .RESET_B(net1001),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_gpio_edge ));
 sky130_fd_sc_hd__dfrtp_1 _11412_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2186),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11413_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2132),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11414_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2177),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11415_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2110),
    .RESET_B(net984),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_hold ));
 sky130_fd_sc_hd__dfrtp_1 _11416_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2138),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11417_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2111),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_mode[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11418_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2130),
    .RESET_B(net984),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_inv ));
 sky130_fd_sc_hd__dfrtp_1 _11419_ (.CLK(clknet_1_1__leaf__04565_),
    .D(net2212),
    .RESET_B(net1001),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_zeropd ));
 sky130_fd_sc_hd__dfrtp_1 _11420_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2115),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.cfg_comp0_center ));
 sky130_fd_sc_hd__dfrtp_1 _11421_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2118),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.cfg_comp1_center ));
 sky130_fd_sc_hd__dfrtp_1 _11422_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2109),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.cfg_comp2_center ));
 sky130_fd_sc_hd__dfrtp_1 _11423_ (.CLK(clknet_1_0__leaf__04565_),
    .D(net2116),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.cfg_comp3_center ));
 sky130_fd_sc_hd__dfrtp_1 _11424_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2142),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11425_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2182),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11426_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2154),
    .RESET_B(net1017),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11427_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2175),
    .RESET_B(net1017),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11428_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2170),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11429_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2205),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11430_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2179),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11431_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2155),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11432_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2150),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11433_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2189),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11434_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2206),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11435_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2141),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11436_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2200),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11437_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2146),
    .RESET_B(net1006),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11438_ (.CLK(clknet_1_0__leaf__04566_),
    .D(net2199),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11439_ (.CLK(clknet_1_1__leaf__04566_),
    .D(net2160),
    .RESET_B(net1006),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_period[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11440_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2108),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11441_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2102),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11442_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2072),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11443_ (.CLK(clknet_2_1__leaf__04567_),
    .D(net2086),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11444_ (.CLK(clknet_2_1__leaf__04567_),
    .D(net2081),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11445_ (.CLK(clknet_2_1__leaf__04567_),
    .D(net2078),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11446_ (.CLK(clknet_2_1__leaf__04567_),
    .D(net2080),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11447_ (.CLK(clknet_2_1__leaf__04567_),
    .D(net2084),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11448_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2067),
    .RESET_B(net1002),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11449_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2079),
    .RESET_B(net1002),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11450_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2071),
    .RESET_B(net1002),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11451_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2069),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[11] ));
 sky130_fd_sc_hd__dfrtp_2 _11452_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2085),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11453_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2087),
    .RESET_B(net1006),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11454_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2073),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11455_ (.CLK(clknet_2_0__leaf__04567_),
    .D(net2070),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11456_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2068),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11457_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2088),
    .RESET_B(net1013),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11458_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2126),
    .RESET_B(net1013),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11459_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2027),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11460_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2096),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11461_ (.CLK(clknet_2_3__leaf__04567_),
    .D(net2076),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11462_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2083),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11463_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2094),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11464_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2041),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11465_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2049),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11466_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2043),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11467_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2055),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11468_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2060),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11469_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2059),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11470_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2047),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11471_ (.CLK(clknet_2_2__leaf__04567_),
    .D(net2040),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11472_ (.CLK(clknet_1_0__leaf__04571_),
    .D(net1428),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11473_ (.CLK(clknet_1_0__leaf__04571_),
    .D(net1421),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11474_ (.CLK(clknet_1_0__leaf__04571_),
    .D(net1289),
    .RESET_B(net981),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11475_ (.CLK(clknet_1_1__leaf__04571_),
    .D(net1646),
    .RESET_B(net982),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11476_ (.CLK(clknet_1_1__leaf__04571_),
    .D(net1639),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11477_ (.CLK(clknet_1_1__leaf__04571_),
    .D(net1631),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11478_ (.CLK(clknet_1_0__leaf__04571_),
    .D(net1624),
    .RESET_B(net982),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11479_ (.CLK(clknet_1_1__leaf__04571_),
    .D(net1616),
    .RESET_B(net982),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11480_ (.CLK(clknet_1_1__leaf__04570_),
    .D(net1300),
    .RESET_B(net1009),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11481_ (.CLK(clknet_1_1__leaf__04570_),
    .D(net1578),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11482_ (.CLK(clknet_1_1__leaf__04570_),
    .D(net1493),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11483_ (.CLK(clknet_1_1__leaf__04570_),
    .D(net1470),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11484_ (.CLK(clknet_1_0__leaf__04570_),
    .D(net1464),
    .RESET_B(net1000),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11485_ (.CLK(clknet_1_0__leaf__04570_),
    .D(net1453),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11486_ (.CLK(clknet_1_0__leaf__04570_),
    .D(net1447),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11487_ (.CLK(clknet_1_0__leaf__04570_),
    .D(net1439),
    .RESET_B(net1001),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11488_ (.CLK(clknet_1_1__leaf__04569_),
    .D(net1540),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11489_ (.CLK(clknet_1_0__leaf__04569_),
    .D(net1533),
    .RESET_B(net979),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11490_ (.CLK(clknet_1_1__leaf__04569_),
    .D(net1525),
    .RESET_B(net989),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11491_ (.CLK(clknet_1_0__leaf__04569_),
    .D(net1518),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11492_ (.CLK(clknet_1_1__leaf__04569_),
    .D(net1511),
    .RESET_B(net989),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11493_ (.CLK(clknet_1_0__leaf__04569_),
    .D(net1504),
    .RESET_B(net989),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11494_ (.CLK(clknet_1_1__leaf__04569_),
    .D(net1487),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11495_ (.CLK(clknet_1_0__leaf__04569_),
    .D(net1480),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11496_ (.CLK(clknet_1_0__leaf__04568_),
    .D(net1607),
    .RESET_B(net987),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11497_ (.CLK(clknet_1_1__leaf__04568_),
    .D(net1600),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11498_ (.CLK(clknet_1_1__leaf__04568_),
    .D(net1591),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11499_ (.CLK(clknet_1_1__leaf__04568_),
    .D(net1583),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11500_ (.CLK(clknet_1_0__leaf__04568_),
    .D(net1568),
    .RESET_B(net987),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11501_ (.CLK(clknet_1_1__leaf__04568_),
    .D(net1561),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11502_ (.CLK(clknet_1_0__leaf__04568_),
    .D(net1553),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11503_ (.CLK(clknet_1_0__leaf__04568_),
    .D(net1546),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11504_ (.CLK(clknet_1_1__leaf__04575_),
    .D(net1432),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11505_ (.CLK(clknet_1_0__leaf__04575_),
    .D(net1421),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11506_ (.CLK(clknet_1_0__leaf__04575_),
    .D(net1289),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11507_ (.CLK(clknet_1_1__leaf__04575_),
    .D(net1646),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11508_ (.CLK(clknet_1_0__leaf__04575_),
    .D(net1641),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11509_ (.CLK(clknet_1_1__leaf__04575_),
    .D(net1635),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11510_ (.CLK(clknet_1_0__leaf__04575_),
    .D(net1624),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11511_ (.CLK(clknet_1_1__leaf__04575_),
    .D(net1618),
    .RESET_B(net987),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11512_ (.CLK(clknet_1_1__leaf__04574_),
    .D(net1300),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11513_ (.CLK(clknet_1_1__leaf__04574_),
    .D(net1578),
    .RESET_B(net1009),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11514_ (.CLK(clknet_1_1__leaf__04574_),
    .D(net1493),
    .RESET_B(net1017),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11515_ (.CLK(clknet_1_1__leaf__04574_),
    .D(net1470),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11516_ (.CLK(clknet_1_0__leaf__04574_),
    .D(net1464),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11517_ (.CLK(clknet_1_0__leaf__04574_),
    .D(net1453),
    .RESET_B(net1009),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11518_ (.CLK(clknet_1_0__leaf__04574_),
    .D(net1447),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11519_ (.CLK(clknet_1_0__leaf__04574_),
    .D(net1439),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11520_ (.CLK(clknet_1_0__leaf__04573_),
    .D(net1540),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11521_ (.CLK(clknet_1_1__leaf__04573_),
    .D(net1532),
    .RESET_B(net991),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11522_ (.CLK(clknet_1_0__leaf__04573_),
    .D(net1525),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11523_ (.CLK(clknet_1_1__leaf__04573_),
    .D(net1518),
    .RESET_B(net991),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11524_ (.CLK(clknet_1_0__leaf__04573_),
    .D(net1511),
    .RESET_B(net991),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11525_ (.CLK(clknet_1_0__leaf__04573_),
    .D(net1504),
    .RESET_B(net991),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11526_ (.CLK(clknet_1_1__leaf__04573_),
    .D(net1487),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11527_ (.CLK(clknet_1_1__leaf__04573_),
    .D(net1480),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11528_ (.CLK(clknet_1_0__leaf__04572_),
    .D(net1607),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11529_ (.CLK(clknet_1_1__leaf__04572_),
    .D(net1600),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11530_ (.CLK(clknet_1_0__leaf__04572_),
    .D(net1591),
    .RESET_B(net985),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11531_ (.CLK(clknet_1_1__leaf__04572_),
    .D(net1583),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11532_ (.CLK(clknet_1_0__leaf__04572_),
    .D(net1568),
    .RESET_B(net979),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11533_ (.CLK(clknet_1_1__leaf__04572_),
    .D(net1561),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11534_ (.CLK(clknet_1_1__leaf__04572_),
    .D(net1553),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11535_ (.CLK(clknet_1_0__leaf__04572_),
    .D(net1546),
    .RESET_B(net987),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11536_ (.CLK(clknet_1_0__leaf__04579_),
    .D(net1428),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11537_ (.CLK(clknet_1_0__leaf__04579_),
    .D(net1421),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11538_ (.CLK(clknet_1_0__leaf__04579_),
    .D(net1289),
    .RESET_B(net999),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11539_ (.CLK(clknet_1_1__leaf__04579_),
    .D(net1646),
    .RESET_B(net1003),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11540_ (.CLK(clknet_1_1__leaf__04579_),
    .D(net1639),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11541_ (.CLK(clknet_1_1__leaf__04579_),
    .D(net1631),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11542_ (.CLK(clknet_1_1__leaf__04579_),
    .D(net1626),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11543_ (.CLK(clknet_1_0__leaf__04579_),
    .D(net1616),
    .RESET_B(net984),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11544_ (.CLK(clknet_1_0__leaf__04578_),
    .D(net1300),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11545_ (.CLK(clknet_1_1__leaf__04578_),
    .D(net1578),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11546_ (.CLK(clknet_1_1__leaf__04578_),
    .D(net1493),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11547_ (.CLK(clknet_1_1__leaf__04578_),
    .D(net1470),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11548_ (.CLK(clknet_1_0__leaf__04578_),
    .D(net1464),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11549_ (.CLK(clknet_1_0__leaf__04578_),
    .D(net1453),
    .RESET_B(net1008),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11550_ (.CLK(clknet_1_0__leaf__04578_),
    .D(net1447),
    .RESET_B(net1004),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11551_ (.CLK(clknet_1_1__leaf__04578_),
    .D(net1439),
    .RESET_B(net1005),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11552_ (.CLK(clknet_1_0__leaf__04577_),
    .D(net1540),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11553_ (.CLK(clknet_1_1__leaf__04577_),
    .D(net1532),
    .RESET_B(net1021),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11554_ (.CLK(clknet_1_0__leaf__04577_),
    .D(net1525),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11555_ (.CLK(clknet_1_1__leaf__04577_),
    .D(net1518),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11556_ (.CLK(clknet_1_0__leaf__04577_),
    .D(net1511),
    .RESET_B(net991),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11557_ (.CLK(clknet_1_0__leaf__04577_),
    .D(net1504),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11558_ (.CLK(clknet_1_1__leaf__04577_),
    .D(net1487),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11559_ (.CLK(clknet_1_1__leaf__04577_),
    .D(net1480),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11560_ (.CLK(clknet_1_0__leaf__04576_),
    .D(net1609),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11561_ (.CLK(clknet_1_0__leaf__04576_),
    .D(net1600),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11562_ (.CLK(clknet_1_0__leaf__04576_),
    .D(net1591),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11563_ (.CLK(clknet_1_1__leaf__04576_),
    .D(net1583),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11564_ (.CLK(clknet_1_0__leaf__04576_),
    .D(net1568),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11565_ (.CLK(clknet_1_1__leaf__04576_),
    .D(net1561),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11566_ (.CLK(clknet_1_1__leaf__04576_),
    .D(net1553),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11567_ (.CLK(clknet_1_1__leaf__04576_),
    .D(net1546),
    .RESET_B(net996),
    .Q(\u_pwm.u_pwm_0.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11568_ (.CLK(clknet_1_1__leaf__04583_),
    .D(net1432),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11569_ (.CLK(clknet_1_0__leaf__04583_),
    .D(net1421),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11570_ (.CLK(clknet_1_0__leaf__04583_),
    .D(net1289),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11571_ (.CLK(clknet_1_0__leaf__04583_),
    .D(net1646),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__dfrtp_2 _11572_ (.CLK(clknet_1_0__leaf__04583_),
    .D(net1639),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11573_ (.CLK(clknet_1_1__leaf__04583_),
    .D(net1631),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11574_ (.CLK(clknet_1_1__leaf__04583_),
    .D(net1626),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11575_ (.CLK(clknet_1_1__leaf__04583_),
    .D(net1618),
    .RESET_B(net986),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11576_ (.CLK(clknet_1_1__leaf__04582_),
    .D(net1301),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11577_ (.CLK(clknet_1_1__leaf__04582_),
    .D(net1578),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11578_ (.CLK(clknet_1_1__leaf__04582_),
    .D(net1493),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11579_ (.CLK(clknet_1_1__leaf__04582_),
    .D(net1470),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11580_ (.CLK(clknet_1_0__leaf__04582_),
    .D(net1464),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11581_ (.CLK(clknet_1_0__leaf__04582_),
    .D(net1453),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11582_ (.CLK(clknet_1_0__leaf__04582_),
    .D(net1447),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11583_ (.CLK(clknet_1_0__leaf__04582_),
    .D(net1439),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11584_ (.CLK(clknet_1_1__leaf__04581_),
    .D(net1540),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11585_ (.CLK(clknet_1_1__leaf__04581_),
    .D(net1532),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11586_ (.CLK(clknet_1_1__leaf__04581_),
    .D(net1525),
    .RESET_B(net990),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11587_ (.CLK(clknet_1_0__leaf__04581_),
    .D(net1518),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11588_ (.CLK(clknet_1_1__leaf__04581_),
    .D(net1511),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11589_ (.CLK(clknet_1_0__leaf__04581_),
    .D(net1504),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[13] ));
 sky130_fd_sc_hd__dfrtp_2 _11590_ (.CLK(clknet_1_0__leaf__04581_),
    .D(net1487),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11591_ (.CLK(clknet_1_0__leaf__04581_),
    .D(net1480),
    .RESET_B(net988),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11592_ (.CLK(clknet_1_0__leaf__04580_),
    .D(net1609),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11593_ (.CLK(clknet_1_0__leaf__04580_),
    .D(net1601),
    .RESET_B(net994),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11594_ (.CLK(clknet_1_0__leaf__04580_),
    .D(net1591),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11595_ (.CLK(clknet_1_1__leaf__04580_),
    .D(net1583),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__dfrtp_2 _11596_ (.CLK(clknet_1_0__leaf__04580_),
    .D(net1568),
    .RESET_B(net993),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11597_ (.CLK(clknet_1_1__leaf__04580_),
    .D(net1561),
    .RESET_B(net995),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11598_ (.CLK(clknet_1_1__leaf__04580_),
    .D(net1554),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11599_ (.CLK(clknet_1_1__leaf__04580_),
    .D(net1546),
    .RESET_B(net997),
    .Q(\u_pwm.u_pwm_0.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11600_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[0] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_pwm0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11601_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[1] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_pwm0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11602_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[2] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_pwm0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11603_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[3] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_pwm0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11604_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[4] ),
    .RESET_B(net1001),
    .Q(\u_pwm.reg_rdata_pwm0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11605_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[5] ),
    .RESET_B(net1007),
    .Q(\u_pwm.reg_rdata_pwm0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11606_ (.CLK(clknet_2_3__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[6] ),
    .RESET_B(net1004),
    .Q(\u_pwm.reg_rdata_pwm0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11607_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[7] ),
    .RESET_B(net1000),
    .Q(\u_pwm.reg_rdata_pwm0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11608_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[8] ),
    .RESET_B(net983),
    .Q(\u_pwm.reg_rdata_pwm0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11609_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[9] ),
    .RESET_B(net983),
    .Q(\u_pwm.reg_rdata_pwm0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11610_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[10] ),
    .RESET_B(net983),
    .Q(\u_pwm.reg_rdata_pwm0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11611_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[11] ),
    .RESET_B(net982),
    .Q(\u_pwm.reg_rdata_pwm0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11612_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[12] ),
    .RESET_B(net982),
    .Q(\u_pwm.reg_rdata_pwm0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11613_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[13] ),
    .RESET_B(net985),
    .Q(\u_pwm.reg_rdata_pwm0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11614_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[14] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11615_ (.CLK(clknet_2_2__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[15] ),
    .RESET_B(net981),
    .Q(\u_pwm.reg_rdata_pwm0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11616_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[16] ),
    .RESET_B(net982),
    .Q(\u_pwm.reg_rdata_pwm0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11617_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[17] ),
    .RESET_B(net985),
    .Q(\u_pwm.reg_rdata_pwm0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11618_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[18] ),
    .RESET_B(net981),
    .Q(\u_pwm.reg_rdata_pwm0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11619_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[19] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11620_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[20] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11621_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[21] ),
    .RESET_B(net980),
    .Q(\u_pwm.reg_rdata_pwm0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11622_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[22] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11623_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[23] ),
    .RESET_B(net980),
    .Q(\u_pwm.reg_rdata_pwm0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11624_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[24] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11625_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[25] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11626_ (.CLK(clknet_2_1__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[26] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11627_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[27] ),
    .RESET_B(net979),
    .Q(\u_pwm.reg_rdata_pwm0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11628_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[28] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11629_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[29] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11630_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[30] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11631_ (.CLK(clknet_2_0__leaf__04564_),
    .D(\u_pwm.u_pwm_0.u_reg.reg_out[31] ),
    .RESET_B(net976),
    .Q(\u_pwm.reg_rdata_pwm0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11632_ (.CLK(clknet_leaf_79_mclk),
    .D(_00352_),
    .RESET_B(net977),
    .Q(\u_pwm.reg_ack_pwm0 ));
 sky130_fd_sc_hd__dfrtp_4 _11633_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00319_),
    .RESET_B(net1016),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11634_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00326_),
    .RESET_B(net1016),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11635_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00327_),
    .RESET_B(net1016),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11636_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00328_),
    .RESET_B(net1040),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11637_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00329_),
    .RESET_B(net1040),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _11638_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00330_),
    .RESET_B(net1040),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11639_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00331_),
    .RESET_B(net1032),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11640_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00332_),
    .RESET_B(net1032),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11641_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00333_),
    .RESET_B(net1032),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11642_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00334_),
    .RESET_B(net1031),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11643_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00320_),
    .RESET_B(net1031),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _11644_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00321_),
    .RESET_B(net1032),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _11645_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00322_),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _11646_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00323_),
    .RESET_B(net1013),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _11647_ (.CLK(clknet_1_0__leaf__04562_),
    .D(_00324_),
    .RESET_B(net1012),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _11648_ (.CLK(clknet_1_1__leaf__04562_),
    .D(_00325_),
    .RESET_B(net1013),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11649_ (.CLK(_04563_),
    .D(\u_pwm.u_pwm_0.u_pwm.pwm_wfm_i ),
    .RESET_B(net983),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_wfm_r ));
 sky130_fd_sc_hd__dfrtp_1 _11650_ (.CLK(clknet_leaf_76_mclk),
    .D(\u_pwm.u_pwm_0.u_pwm.pwm_ovflow ),
    .RESET_B(net1000),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_ovflow_l ));
 sky130_fd_sc_hd__dfrtp_1 _11651_ (.CLK(clknet_leaf_76_mclk),
    .D(_00318_),
    .RESET_B(net1000),
    .Q(\u_pwm.u_pwm_0.gpio_tgr ));
 sky130_fd_sc_hd__dfrtp_1 _11652_ (.CLK(clknet_leaf_76_mclk),
    .D(_00317_),
    .RESET_B(net1000),
    .Q(\u_pwm.u_pwm_0.u_pwm.gpio_l ));
 sky130_fd_sc_hd__dfrtp_1 _11653_ (.CLK(clknet_leaf_73_mclk),
    .D(_00335_),
    .RESET_B(net1010),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11654_ (.CLK(clknet_leaf_74_mclk),
    .D(_00341_),
    .RESET_B(net1010),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11655_ (.CLK(clknet_leaf_74_mclk),
    .D(_00342_),
    .RESET_B(net1010),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11656_ (.CLK(clknet_leaf_73_mclk),
    .D(_00343_),
    .RESET_B(net1010),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11657_ (.CLK(clknet_leaf_73_mclk),
    .D(_00344_),
    .RESET_B(net1010),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11658_ (.CLK(clknet_leaf_73_mclk),
    .D(_00345_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11659_ (.CLK(clknet_leaf_73_mclk),
    .D(_00346_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11660_ (.CLK(clknet_leaf_73_mclk),
    .D(_00347_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11661_ (.CLK(clknet_leaf_73_mclk),
    .D(_00348_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11662_ (.CLK(clknet_leaf_73_mclk),
    .D(_00349_),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11663_ (.CLK(clknet_leaf_72_mclk),
    .D(_00336_),
    .RESET_B(net1014),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11664_ (.CLK(clknet_leaf_72_mclk),
    .D(_00337_),
    .RESET_B(net1016),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11665_ (.CLK(clknet_leaf_72_mclk),
    .D(_00338_),
    .RESET_B(net1016),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11666_ (.CLK(clknet_leaf_72_mclk),
    .D(_00339_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11667_ (.CLK(clknet_leaf_73_mclk),
    .D(_00340_),
    .RESET_B(net1015),
    .Q(\u_pwm.u_pwm_0.u_pwm.pwm_scnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11668_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2125),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_scale[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11669_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2128),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_scale[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11670_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2134),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_scale[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11671_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2123),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_scale[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11672_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2153),
    .RESET_B(net888),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_oneshot ));
 sky130_fd_sc_hd__dfrtp_1 _11673_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2103),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_gpio_enb ));
 sky130_fd_sc_hd__dfrtp_1 _11674_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2137),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_gpio_edge ));
 sky130_fd_sc_hd__dfrtp_1 _11675_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2183),
    .RESET_B(net875),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11676_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2147),
    .RESET_B(net876),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11677_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2201),
    .RESET_B(net875),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11678_ (.CLK(clknet_1_1__leaf__04587_),
    .D(net2140),
    .RESET_B(net874),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_hold ));
 sky130_fd_sc_hd__dfrtp_1 _11679_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2172),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11680_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2217),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11681_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2181),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_inv ));
 sky130_fd_sc_hd__dfrtp_1 _11682_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2207),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_zeropd ));
 sky130_fd_sc_hd__dfrtp_1 _11683_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2124),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_comp0_center ));
 sky130_fd_sc_hd__dfrtp_1 _11684_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2194),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.cfg_comp1_center ));
 sky130_fd_sc_hd__dfrtp_1 _11685_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2204),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_comp2_center ));
 sky130_fd_sc_hd__dfrtp_1 _11686_ (.CLK(clknet_1_0__leaf__04587_),
    .D(net2092),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_comp3_center ));
 sky130_fd_sc_hd__dfrtp_1 _11687_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2254),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11688_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2289),
    .RESET_B(net881),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11689_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2164),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11690_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2233),
    .RESET_B(net881),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11691_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2232),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11692_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2224),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11693_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2215),
    .RESET_B(net885),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11694_ (.CLK(clknet_1_1__leaf__04588_),
    .D(net2241),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11695_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2312),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11696_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2230),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11697_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2275),
    .RESET_B(net886),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11698_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2240),
    .RESET_B(net886),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11699_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2321),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11700_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2272),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11701_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2325),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11702_ (.CLK(clknet_1_0__leaf__04588_),
    .D(net2245),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_period[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11703_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2106),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11704_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2107),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11705_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2101),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11706_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2135),
    .RESET_B(net881),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11707_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2136),
    .RESET_B(net881),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11708_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2093),
    .RESET_B(net893),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11709_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2100),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11710_ (.CLK(clknet_2_3__leaf__04589_),
    .D(net2095),
    .RESET_B(net885),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11711_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2180),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11712_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2178),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__dfrtp_2 _11713_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2145),
    .RESET_B(net889),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11714_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2149),
    .RESET_B(net886),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11715_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2159),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11716_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2176),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[13] ));
 sky130_fd_sc_hd__dfrtp_2 _11717_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2163),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[14] ));
 sky130_fd_sc_hd__dfrtp_2 _11718_ (.CLK(clknet_2_2__leaf__04589_),
    .D(net2119),
    .RESET_B(net883),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11719_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1974),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11720_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1989),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11721_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1975),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11722_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1964),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11723_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net1971),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11724_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1973),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11725_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1972),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11726_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net1987),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11727_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net2075),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11728_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2121),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11729_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2127),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11730_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2113),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11731_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2074),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11732_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2105),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11733_ (.CLK(clknet_2_1__leaf__04589_),
    .D(net2082),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11734_ (.CLK(clknet_2_0__leaf__04589_),
    .D(net2104),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11735_ (.CLK(clknet_1_1__leaf__04593_),
    .D(net1428),
    .RESET_B(net874),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11736_ (.CLK(clknet_1_1__leaf__04593_),
    .D(net1422),
    .RESET_B(net875),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11737_ (.CLK(clknet_1_1__leaf__04593_),
    .D(net1290),
    .RESET_B(net875),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11738_ (.CLK(clknet_1_1__leaf__04593_),
    .D(net1646),
    .RESET_B(net874),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11739_ (.CLK(clknet_1_0__leaf__04593_),
    .D(net1639),
    .RESET_B(net874),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11740_ (.CLK(clknet_1_0__leaf__04593_),
    .D(net1631),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11741_ (.CLK(clknet_1_0__leaf__04593_),
    .D(net1624),
    .RESET_B(net874),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11742_ (.CLK(clknet_1_0__leaf__04593_),
    .D(net1616),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11743_ (.CLK(clknet_1_1__leaf__04592_),
    .D(net1297),
    .RESET_B(net893),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11744_ (.CLK(clknet_1_1__leaf__04592_),
    .D(net1574),
    .RESET_B(net893),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11745_ (.CLK(clknet_1_1__leaf__04592_),
    .D(net1491),
    .RESET_B(net893),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11746_ (.CLK(clknet_1_1__leaf__04592_),
    .D(net1468),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11747_ (.CLK(clknet_1_0__leaf__04592_),
    .D(net1461),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11748_ (.CLK(clknet_1_0__leaf__04592_),
    .D(net1450),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11749_ (.CLK(clknet_1_0__leaf__04592_),
    .D(net1444),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11750_ (.CLK(clknet_1_0__leaf__04592_),
    .D(net1440),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11751_ (.CLK(clknet_1_1__leaf__04591_),
    .D(net1538),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11752_ (.CLK(clknet_1_0__leaf__04591_),
    .D(net1530),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11753_ (.CLK(clknet_1_0__leaf__04591_),
    .D(net1523),
    .RESET_B(net854),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11754_ (.CLK(clknet_1_0__leaf__04591_),
    .D(net1516),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11755_ (.CLK(clknet_1_0__leaf__04591_),
    .D(net1508),
    .RESET_B(net854),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11756_ (.CLK(clknet_1_1__leaf__04591_),
    .D(net1500),
    .RESET_B(net856),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11757_ (.CLK(clknet_1_1__leaf__04591_),
    .D(net1484),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11758_ (.CLK(clknet_1_1__leaf__04591_),
    .D(net1478),
    .RESET_B(net856),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11759_ (.CLK(clknet_1_1__leaf__04590_),
    .D(net1605),
    .RESET_B(net862),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11760_ (.CLK(clknet_1_0__leaf__04590_),
    .D(net1596),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11761_ (.CLK(clknet_1_1__leaf__04590_),
    .D(net1588),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11762_ (.CLK(clknet_1_0__leaf__04590_),
    .D(net1580),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11763_ (.CLK(clknet_1_1__leaf__04590_),
    .D(net1564),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11764_ (.CLK(clknet_1_1__leaf__04590_),
    .D(net1558),
    .RESET_B(net860),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11765_ (.CLK(clknet_1_0__leaf__04590_),
    .D(net1551),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11766_ (.CLK(clknet_1_0__leaf__04590_),
    .D(net1544),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11767_ (.CLK(clknet_1_1__leaf__04597_),
    .D(net1428),
    .RESET_B(net873),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11768_ (.CLK(clknet_1_1__leaf__04597_),
    .D(net1422),
    .RESET_B(net873),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11769_ (.CLK(clknet_1_1__leaf__04597_),
    .D(net1290),
    .RESET_B(net876),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11770_ (.CLK(clknet_1_1__leaf__04597_),
    .D(net1648),
    .RESET_B(net873),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11771_ (.CLK(clknet_1_0__leaf__04597_),
    .D(net1639),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11772_ (.CLK(clknet_1_0__leaf__04597_),
    .D(net1631),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11773_ (.CLK(clknet_1_0__leaf__04597_),
    .D(net1624),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11774_ (.CLK(clknet_1_0__leaf__04597_),
    .D(net1616),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11775_ (.CLK(clknet_1_1__leaf__04596_),
    .D(net1297),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11776_ (.CLK(clknet_1_1__leaf__04596_),
    .D(net1574),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11777_ (.CLK(clknet_1_1__leaf__04596_),
    .D(net1491),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11778_ (.CLK(clknet_1_1__leaf__04596_),
    .D(net1468),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11779_ (.CLK(clknet_1_0__leaf__04596_),
    .D(net1460),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11780_ (.CLK(clknet_1_0__leaf__04596_),
    .D(net1451),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11781_ (.CLK(clknet_1_0__leaf__04596_),
    .D(net1444),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11782_ (.CLK(clknet_1_0__leaf__04596_),
    .D(net1436),
    .RESET_B(net885),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11783_ (.CLK(clknet_1_1__leaf__04595_),
    .D(net1538),
    .RESET_B(net856),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11784_ (.CLK(clknet_1_0__leaf__04595_),
    .D(net1530),
    .RESET_B(net854),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11785_ (.CLK(clknet_1_0__leaf__04595_),
    .D(net1523),
    .RESET_B(net854),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11786_ (.CLK(clknet_1_0__leaf__04595_),
    .D(net1515),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11787_ (.CLK(clknet_1_0__leaf__04595_),
    .D(net1508),
    .RESET_B(net860),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11788_ (.CLK(clknet_1_1__leaf__04595_),
    .D(net1500),
    .RESET_B(net856),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11789_ (.CLK(clknet_1_1__leaf__04595_),
    .D(net1484),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11790_ (.CLK(clknet_1_1__leaf__04595_),
    .D(net1478),
    .RESET_B(net865),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11791_ (.CLK(clknet_1_1__leaf__04594_),
    .D(net1605),
    .RESET_B(net834),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11792_ (.CLK(clknet_1_0__leaf__04594_),
    .D(net1596),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11793_ (.CLK(clknet_1_1__leaf__04594_),
    .D(net1588),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11794_ (.CLK(clknet_1_0__leaf__04594_),
    .D(net1580),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11795_ (.CLK(clknet_1_1__leaf__04594_),
    .D(net1565),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11796_ (.CLK(clknet_1_0__leaf__04594_),
    .D(net1558),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11797_ (.CLK(clknet_1_0__leaf__04594_),
    .D(net1551),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11798_ (.CLK(clknet_1_1__leaf__04594_),
    .D(net1544),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11799_ (.CLK(clknet_1_1__leaf__04601_),
    .D(net1432),
    .RESET_B(net876),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11800_ (.CLK(clknet_1_1__leaf__04601_),
    .D(net1422),
    .RESET_B(net876),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11801_ (.CLK(clknet_1_1__leaf__04601_),
    .D(net1290),
    .RESET_B(net876),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11802_ (.CLK(clknet_1_1__leaf__04601_),
    .D(net1648),
    .RESET_B(net873),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11803_ (.CLK(clknet_1_0__leaf__04601_),
    .D(net1641),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11804_ (.CLK(clknet_1_0__leaf__04601_),
    .D(net1635),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11805_ (.CLK(clknet_1_0__leaf__04601_),
    .D(net1624),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11806_ (.CLK(clknet_1_0__leaf__04601_),
    .D(net1616),
    .RESET_B(net872),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11807_ (.CLK(clknet_1_1__leaf__04600_),
    .D(net1297),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11808_ (.CLK(clknet_1_0__leaf__04600_),
    .D(net1575),
    .RESET_B(net891),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11809_ (.CLK(clknet_1_0__leaf__04600_),
    .D(net1491),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11810_ (.CLK(clknet_1_0__leaf__04600_),
    .D(net1469),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11811_ (.CLK(clknet_1_0__leaf__04600_),
    .D(net1460),
    .RESET_B(net890),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11812_ (.CLK(clknet_1_1__leaf__04600_),
    .D(net1451),
    .RESET_B(net893),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11813_ (.CLK(clknet_1_1__leaf__04600_),
    .D(net1445),
    .RESET_B(net887),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11814_ (.CLK(clknet_1_1__leaf__04600_),
    .D(net1440),
    .RESET_B(net885),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11815_ (.CLK(clknet_1_0__leaf__04599_),
    .D(net1537),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11816_ (.CLK(clknet_1_0__leaf__04599_),
    .D(net1529),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11817_ (.CLK(clknet_1_1__leaf__04599_),
    .D(net1522),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11818_ (.CLK(clknet_1_0__leaf__04599_),
    .D(net1515),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11819_ (.CLK(clknet_1_1__leaf__04599_),
    .D(net1508),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11820_ (.CLK(clknet_1_1__leaf__04599_),
    .D(net1500),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11821_ (.CLK(clknet_1_1__leaf__04599_),
    .D(net1484),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11822_ (.CLK(clknet_1_0__leaf__04599_),
    .D(net1477),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11823_ (.CLK(clknet_1_1__leaf__04598_),
    .D(net1605),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11824_ (.CLK(clknet_1_0__leaf__04598_),
    .D(net1597),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11825_ (.CLK(clknet_1_1__leaf__04598_),
    .D(net1588),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11826_ (.CLK(clknet_1_0__leaf__04598_),
    .D(net1580),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11827_ (.CLK(clknet_1_1__leaf__04598_),
    .D(net1565),
    .RESET_B(net834),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11828_ (.CLK(clknet_1_0__leaf__04598_),
    .D(net1558),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11829_ (.CLK(clknet_1_0__leaf__04598_),
    .D(net1551),
    .RESET_B(net833),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11830_ (.CLK(clknet_1_1__leaf__04598_),
    .D(net1544),
    .RESET_B(net834),
    .Q(\u_pwm.u_pwm_1.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11831_ (.CLK(clknet_1_1__leaf__04605_),
    .D(net1428),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__dfrtp_2 _11832_ (.CLK(clknet_1_0__leaf__04605_),
    .D(net1421),
    .RESET_B(net865),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11833_ (.CLK(clknet_1_1__leaf__04605_),
    .D(net1289),
    .RESET_B(net882),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11834_ (.CLK(clknet_1_1__leaf__04605_),
    .D(net1646),
    .RESET_B(net882),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11835_ (.CLK(clknet_1_0__leaf__04605_),
    .D(net1639),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[12] ));
 sky130_fd_sc_hd__dfrtp_2 _11836_ (.CLK(clknet_1_0__leaf__04605_),
    .D(net1631),
    .RESET_B(net865),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11837_ (.CLK(clknet_1_1__leaf__04605_),
    .D(net1624),
    .RESET_B(net865),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11838_ (.CLK(clknet_1_0__leaf__04605_),
    .D(net1613),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11839_ (.CLK(clknet_1_1__leaf__04604_),
    .D(net1297),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11840_ (.CLK(clknet_1_0__leaf__04604_),
    .D(net1574),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11841_ (.CLK(clknet_1_1__leaf__04604_),
    .D(net1491),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11842_ (.CLK(clknet_1_0__leaf__04604_),
    .D(net1469),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11843_ (.CLK(clknet_1_0__leaf__04604_),
    .D(net1460),
    .RESET_B(net879),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11844_ (.CLK(clknet_1_0__leaf__04604_),
    .D(net1451),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11845_ (.CLK(clknet_1_1__leaf__04604_),
    .D(net1445),
    .RESET_B(net885),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11846_ (.CLK(clknet_1_1__leaf__04604_),
    .D(net1436),
    .RESET_B(net884),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__dfrtp_2 _11847_ (.CLK(clknet_1_1__leaf__04603_),
    .D(net1538),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11848_ (.CLK(clknet_1_1__leaf__04603_),
    .D(net1530),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11849_ (.CLK(clknet_1_1__leaf__04603_),
    .D(net1523),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__dfrtp_2 _11850_ (.CLK(clknet_1_0__leaf__04603_),
    .D(net1516),
    .RESET_B(net860),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11851_ (.CLK(clknet_1_0__leaf__04603_),
    .D(net1508),
    .RESET_B(net860),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11852_ (.CLK(clknet_1_0__leaf__04603_),
    .D(net1500),
    .RESET_B(net860),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11853_ (.CLK(clknet_1_0__leaf__04603_),
    .D(net1484),
    .RESET_B(net859),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[14] ));
 sky130_fd_sc_hd__dfrtp_2 _11854_ (.CLK(clknet_1_1__leaf__04603_),
    .D(net1479),
    .RESET_B(net863),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__dfrtp_2 _11855_ (.CLK(clknet_1_0__leaf__04602_),
    .D(net1605),
    .RESET_B(net862),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__dfrtp_2 _11856_ (.CLK(clknet_1_0__leaf__04602_),
    .D(net1597),
    .RESET_B(net862),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11857_ (.CLK(clknet_1_1__leaf__04602_),
    .D(net1588),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__dfrtp_2 _11858_ (.CLK(clknet_1_0__leaf__04602_),
    .D(net1580),
    .RESET_B(net862),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11859_ (.CLK(clknet_1_1__leaf__04602_),
    .D(net1565),
    .RESET_B(net864),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11860_ (.CLK(clknet_1_1__leaf__04602_),
    .D(net1558),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11861_ (.CLK(clknet_1_1__leaf__04602_),
    .D(net1551),
    .RESET_B(net861),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11862_ (.CLK(clknet_1_0__leaf__04602_),
    .D(net1544),
    .RESET_B(net862),
    .Q(\u_pwm.u_pwm_1.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11863_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[0] ),
    .RESET_B(net895),
    .Q(\u_pwm.reg_rdata_pwm1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11864_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[1] ),
    .RESET_B(net893),
    .Q(\u_pwm.reg_rdata_pwm1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11865_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[2] ),
    .RESET_B(net893),
    .Q(\u_pwm.reg_rdata_pwm1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11866_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[3] ),
    .RESET_B(net895),
    .Q(\u_pwm.reg_rdata_pwm1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11867_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[4] ),
    .RESET_B(net884),
    .Q(\u_pwm.reg_rdata_pwm1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11868_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[5] ),
    .RESET_B(net888),
    .Q(\u_pwm.reg_rdata_pwm1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11869_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[6] ),
    .RESET_B(net887),
    .Q(\u_pwm.reg_rdata_pwm1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11870_ (.CLK(clknet_2_3__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[7] ),
    .RESET_B(net887),
    .Q(\u_pwm.reg_rdata_pwm1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11871_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[8] ),
    .RESET_B(net873),
    .Q(\u_pwm.reg_rdata_pwm1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11872_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[9] ),
    .RESET_B(net876),
    .Q(\u_pwm.reg_rdata_pwm1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11873_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[10] ),
    .RESET_B(net876),
    .Q(\u_pwm.reg_rdata_pwm1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11874_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[11] ),
    .RESET_B(net874),
    .Q(\u_pwm.reg_rdata_pwm1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11875_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[12] ),
    .RESET_B(net874),
    .Q(\u_pwm.reg_rdata_pwm1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11876_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[13] ),
    .RESET_B(net874),
    .Q(\u_pwm.reg_rdata_pwm1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11877_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[14] ),
    .RESET_B(net874),
    .Q(\u_pwm.reg_rdata_pwm1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11878_ (.CLK(clknet_2_2__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[15] ),
    .RESET_B(net874),
    .Q(\u_pwm.reg_rdata_pwm1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11879_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[16] ),
    .RESET_B(net862),
    .Q(\u_pwm.reg_rdata_pwm1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _11880_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[17] ),
    .RESET_B(net859),
    .Q(\u_pwm.reg_rdata_pwm1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _11881_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[18] ),
    .RESET_B(net864),
    .Q(\u_pwm.reg_rdata_pwm1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _11882_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[19] ),
    .RESET_B(net861),
    .Q(\u_pwm.reg_rdata_pwm1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _11883_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[20] ),
    .RESET_B(net863),
    .Q(\u_pwm.reg_rdata_pwm1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _11884_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[21] ),
    .RESET_B(net860),
    .Q(\u_pwm.reg_rdata_pwm1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _11885_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[22] ),
    .RESET_B(net859),
    .Q(\u_pwm.reg_rdata_pwm1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _11886_ (.CLK(clknet_2_1__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[23] ),
    .RESET_B(net859),
    .Q(\u_pwm.reg_rdata_pwm1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _11887_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[24] ),
    .RESET_B(net855),
    .Q(\u_pwm.reg_rdata_pwm1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _11888_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[25] ),
    .RESET_B(net854),
    .Q(\u_pwm.reg_rdata_pwm1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _11889_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[26] ),
    .RESET_B(net852),
    .Q(\u_pwm.reg_rdata_pwm1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _11890_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[27] ),
    .RESET_B(net855),
    .Q(\u_pwm.reg_rdata_pwm1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _11891_ (.CLK(clknet_2_0__leaf__04586_),
    .D(net2203),
    .RESET_B(net855),
    .Q(\u_pwm.reg_rdata_pwm1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _11892_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[29] ),
    .RESET_B(net857),
    .Q(\u_pwm.reg_rdata_pwm1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _11893_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[30] ),
    .RESET_B(net852),
    .Q(\u_pwm.reg_rdata_pwm1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _11894_ (.CLK(clknet_2_0__leaf__04586_),
    .D(\u_pwm.u_pwm_1.u_reg.reg_out[31] ),
    .RESET_B(net856),
    .Q(\u_pwm.reg_rdata_pwm1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _11895_ (.CLK(clknet_leaf_80_mclk),
    .D(_00405_),
    .RESET_B(net977),
    .Q(\u_pwm.reg_ack_pwm1 ));
 sky130_fd_sc_hd__dfrtp_4 _11896_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00372_),
    .RESET_B(net880),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _11897_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00379_),
    .RESET_B(net880),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _11898_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00380_),
    .RESET_B(net880),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _11899_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00381_),
    .RESET_B(net880),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _11900_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00382_),
    .RESET_B(net850),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11901_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00383_),
    .RESET_B(net850),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _11902_ (.CLK(clknet_1_1__leaf__04584_),
    .D(_00384_),
    .RESET_B(net850),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _11903_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00385_),
    .RESET_B(net849),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _11904_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00386_),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _11905_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00387_),
    .RESET_B(net846),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_4 _11906_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00373_),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _11907_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00374_),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _11908_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00375_),
    .RESET_B(net846),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _11909_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00376_),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_4 _11910_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00377_),
    .RESET_B(net847),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_4 _11911_ (.CLK(clknet_1_0__leaf__04584_),
    .D(_00378_),
    .RESET_B(net848),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11912_ (.CLK(_04585_),
    .D(\u_pwm.u_pwm_1.u_pwm.pwm_wfm_i ),
    .RESET_B(net865),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_wfm_r ));
 sky130_fd_sc_hd__dfrtp_1 _11913_ (.CLK(clknet_leaf_86_mclk),
    .D(\u_pwm.u_pwm_1.u_pwm.pwm_ovflow ),
    .RESET_B(net889),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_ovflow_l ));
 sky130_fd_sc_hd__dfrtp_1 _11914_ (.CLK(clknet_leaf_87_mclk),
    .D(_00371_),
    .RESET_B(net889),
    .Q(\u_pwm.u_pwm_1.gpio_tgr ));
 sky130_fd_sc_hd__dfrtp_1 _11915_ (.CLK(clknet_leaf_87_mclk),
    .D(_00370_),
    .RESET_B(net889),
    .Q(\u_pwm.u_pwm_1.u_pwm.gpio_l ));
 sky130_fd_sc_hd__dfrtp_1 _11916_ (.CLK(clknet_leaf_88_mclk),
    .D(_00388_),
    .RESET_B(net895),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11917_ (.CLK(clknet_leaf_89_mclk),
    .D(_00394_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11918_ (.CLK(clknet_leaf_89_mclk),
    .D(_00395_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11919_ (.CLK(clknet_leaf_88_mclk),
    .D(_00396_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11920_ (.CLK(clknet_leaf_88_mclk),
    .D(_00397_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11921_ (.CLK(clknet_leaf_88_mclk),
    .D(_00398_),
    .RESET_B(net895),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11922_ (.CLK(clknet_leaf_88_mclk),
    .D(_00399_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11923_ (.CLK(clknet_leaf_89_mclk),
    .D(_00400_),
    .RESET_B(net894),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11924_ (.CLK(clknet_leaf_90_mclk),
    .D(_00401_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11925_ (.CLK(clknet_leaf_90_mclk),
    .D(_00402_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11926_ (.CLK(clknet_leaf_90_mclk),
    .D(_00389_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11927_ (.CLK(clknet_leaf_89_mclk),
    .D(_00390_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11928_ (.CLK(clknet_leaf_89_mclk),
    .D(_00391_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11929_ (.CLK(clknet_leaf_89_mclk),
    .D(_00392_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11930_ (.CLK(clknet_leaf_89_mclk),
    .D(_00393_),
    .RESET_B(net892),
    .Q(\u_pwm.u_pwm_1.u_pwm.pwm_scnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11931_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2211),
    .RESET_B(net842),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_scale[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11932_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2220),
    .RESET_B(net842),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_scale[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11933_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2221),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_scale[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11934_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2218),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_scale[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11935_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2229),
    .RESET_B(net844),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_oneshot ));
 sky130_fd_sc_hd__dfrtp_1 _11936_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2219),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_gpio_enb ));
 sky130_fd_sc_hd__dfrtp_1 _11937_ (.CLK(clknet_1_1__leaf__04609_),
    .D(net2225),
    .RESET_B(net844),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_gpio_edge ));
 sky130_fd_sc_hd__dfrtp_4 _11938_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[8] ),
    .RESET_B(net832),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11939_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[9] ),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[1] ));
 sky130_fd_sc_hd__dfrtp_2 _11940_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[10] ),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_gpio_sel[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11941_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[11] ),
    .RESET_B(net853),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_hold ));
 sky130_fd_sc_hd__dfrtp_1 _11942_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[12] ),
    .RESET_B(net823),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_mode[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11943_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[13] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11944_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[14] ),
    .RESET_B(net852),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_inv ));
 sky130_fd_sc_hd__dfrtp_1 _11945_ (.CLK(clknet_1_0__leaf__04609_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_0[15] ),
    .RESET_B(net825),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_zeropd ));
 sky130_fd_sc_hd__dfrtp_1 _11946_ (.CLK(clknet_1_0__leaf__04609_),
    .D(net2235),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.cfg_comp0_center ));
 sky130_fd_sc_hd__dfrtp_1 _11947_ (.CLK(clknet_1_0__leaf__04609_),
    .D(net2262),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_comp1_center ));
 sky130_fd_sc_hd__dfrtp_1 _11948_ (.CLK(clknet_1_0__leaf__04609_),
    .D(net2234),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_comp2_center ));
 sky130_fd_sc_hd__dfrtp_1 _11949_ (.CLK(clknet_1_0__leaf__04609_),
    .D(net2339),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_comp3_center ));
 sky130_fd_sc_hd__dfrtp_1 _11950_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2151),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11951_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2139),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11952_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2143),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11953_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2148),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11954_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2152),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11955_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2162),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11956_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2185),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11957_ (.CLK(clknet_1_1__leaf__04610_),
    .D(net2173),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11958_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[8] ),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11959_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[9] ),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11960_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[10] ),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11961_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[11] ),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11962_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[12] ),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11963_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[13] ),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11964_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[14] ),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11965_ (.CLK(clknet_1_0__leaf__04610_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_1[15] ),
    .RESET_B(net817),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_period[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11966_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2197),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11967_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2208),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11968_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2196),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11969_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2222),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11970_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2227),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[4] ));
 sky130_fd_sc_hd__dfrtp_2 _11971_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2129),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[5] ));
 sky130_fd_sc_hd__dfrtp_2 _11972_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2117),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[6] ));
 sky130_fd_sc_hd__dfrtp_2 _11973_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2131),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11974_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[8] ),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11975_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[9] ),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11976_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[10] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11977_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[11] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11978_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[12] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11979_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[13] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11980_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[14] ),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11981_ (.CLK(clknet_2_1__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[15] ),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11982_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2161),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _11983_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2169),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _11984_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2210),
    .RESET_B(net821),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _11985_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2209),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _11986_ (.CLK(clknet_2_3__leaf__04611_),
    .D(net2216),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _11987_ (.CLK(clknet_2_2__leaf__04611_),
    .D(net2334),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _11988_ (.CLK(clknet_2_0__leaf__04611_),
    .D(net2276),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _11989_ (.CLK(clknet_2_0__leaf__04611_),
    .D(net2213),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _11990_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[24] ),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11991_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[25] ),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _11992_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[26] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _11993_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[27] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _11994_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[28] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _11995_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[29] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _11996_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[30] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _11997_ (.CLK(clknet_2_0__leaf__04611_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_2[31] ),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _11998_ (.CLK(clknet_1_0__leaf__04615_),
    .D(net1428),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[8] ));
 sky130_fd_sc_hd__dfrtp_1 _11999_ (.CLK(clknet_1_1__leaf__04615_),
    .D(net1421),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12000_ (.CLK(clknet_1_1__leaf__04615_),
    .D(net1289),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12001_ (.CLK(clknet_1_1__leaf__04615_),
    .D(net1646),
    .RESET_B(net852),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12002_ (.CLK(clknet_1_0__leaf__04615_),
    .D(net1639),
    .RESET_B(net823),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12003_ (.CLK(clknet_1_0__leaf__04615_),
    .D(net1631),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12004_ (.CLK(clknet_1_1__leaf__04615_),
    .D(net1624),
    .RESET_B(net852),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12005_ (.CLK(clknet_1_0__leaf__04615_),
    .D(net1613),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12006_ (.CLK(clknet_1_0__leaf__04614_),
    .D(net1295),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12007_ (.CLK(clknet_1_0__leaf__04614_),
    .D(net1573),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12008_ (.CLK(clknet_1_0__leaf__04614_),
    .D(net1492),
    .RESET_B(net842),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12009_ (.CLK(clknet_1_0__leaf__04614_),
    .D(net1468),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12010_ (.CLK(clknet_1_1__leaf__04614_),
    .D(net1459),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12011_ (.CLK(clknet_1_1__leaf__04614_),
    .D(net1451),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12012_ (.CLK(clknet_1_1__leaf__04614_),
    .D(net1443),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12013_ (.CLK(clknet_1_1__leaf__04614_),
    .D(net1435),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12014_ (.CLK(clknet_1_1__leaf__04613_),
    .D(net1536),
    .RESET_B(net767),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12015_ (.CLK(clknet_1_0__leaf__04613_),
    .D(net1528),
    .RESET_B(net761),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12016_ (.CLK(clknet_1_0__leaf__04613_),
    .D(net1521),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12017_ (.CLK(clknet_1_1__leaf__04613_),
    .D(net1514),
    .RESET_B(net767),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12018_ (.CLK(clknet_1_1__leaf__04613_),
    .D(net1507),
    .RESET_B(net768),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12019_ (.CLK(clknet_1_0__leaf__04613_),
    .D(net1502),
    .RESET_B(net761),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12020_ (.CLK(clknet_1_0__leaf__04613_),
    .D(net1483),
    .RESET_B(net767),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12021_ (.CLK(clknet_1_1__leaf__04613_),
    .D(net1476),
    .RESET_B(net767),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12022_ (.CLK(clknet_1_0__leaf__04612_),
    .D(net1605),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12023_ (.CLK(clknet_1_0__leaf__04612_),
    .D(net1597),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12024_ (.CLK(clknet_1_0__leaf__04612_),
    .D(net1588),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12025_ (.CLK(clknet_1_0__leaf__04612_),
    .D(net1580),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12026_ (.CLK(clknet_1_1__leaf__04612_),
    .D(net1565),
    .RESET_B(net830),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12027_ (.CLK(clknet_1_1__leaf__04612_),
    .D(net1558),
    .RESET_B(net832),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12028_ (.CLK(clknet_1_1__leaf__04612_),
    .D(net1551),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12029_ (.CLK(clknet_1_1__leaf__04612_),
    .D(net1544),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_0[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12030_ (.CLK(clknet_1_1__leaf__04619_),
    .D(net1428),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12031_ (.CLK(clknet_1_1__leaf__04619_),
    .D(net1421),
    .RESET_B(net827),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12032_ (.CLK(clknet_1_0__leaf__04619_),
    .D(net1289),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12033_ (.CLK(clknet_1_1__leaf__04619_),
    .D(net1646),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12034_ (.CLK(clknet_1_0__leaf__04619_),
    .D(net1639),
    .RESET_B(net825),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12035_ (.CLK(clknet_1_0__leaf__04619_),
    .D(net1631),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12036_ (.CLK(clknet_1_1__leaf__04619_),
    .D(net1624),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12037_ (.CLK(clknet_1_0__leaf__04619_),
    .D(net1617),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12038_ (.CLK(clknet_1_1__leaf__04618_),
    .D(net1295),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12039_ (.CLK(clknet_1_1__leaf__04618_),
    .D(net1573),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12040_ (.CLK(clknet_1_1__leaf__04618_),
    .D(net1492),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12041_ (.CLK(clknet_1_0__leaf__04618_),
    .D(net1468),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12042_ (.CLK(clknet_1_0__leaf__04618_),
    .D(net1459),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12043_ (.CLK(clknet_1_1__leaf__04618_),
    .D(net1451),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12044_ (.CLK(clknet_1_0__leaf__04618_),
    .D(net1443),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12045_ (.CLK(clknet_1_0__leaf__04618_),
    .D(net1435),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12046_ (.CLK(clknet_1_1__leaf__04617_),
    .D(net1536),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12047_ (.CLK(clknet_1_0__leaf__04617_),
    .D(net1528),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12048_ (.CLK(clknet_1_0__leaf__04617_),
    .D(net1521),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12049_ (.CLK(clknet_1_0__leaf__04617_),
    .D(net1514),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12050_ (.CLK(clknet_1_1__leaf__04617_),
    .D(net1507),
    .RESET_B(net761),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12051_ (.CLK(clknet_1_1__leaf__04617_),
    .D(net1502),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12052_ (.CLK(clknet_1_0__leaf__04617_),
    .D(net1483),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12053_ (.CLK(clknet_1_1__leaf__04617_),
    .D(net1476),
    .RESET_B(net761),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12054_ (.CLK(clknet_1_0__leaf__04616_),
    .D(net1605),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12055_ (.CLK(clknet_1_0__leaf__04616_),
    .D(net1597),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12056_ (.CLK(clknet_1_0__leaf__04616_),
    .D(net1588),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12057_ (.CLK(clknet_1_1__leaf__04616_),
    .D(net1580),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12058_ (.CLK(clknet_1_1__leaf__04616_),
    .D(net1565),
    .RESET_B(net830),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12059_ (.CLK(clknet_1_1__leaf__04616_),
    .D(net1558),
    .RESET_B(net832),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12060_ (.CLK(clknet_1_1__leaf__04616_),
    .D(net1551),
    .RESET_B(net832),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12061_ (.CLK(clknet_1_0__leaf__04616_),
    .D(net1544),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_1[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12062_ (.CLK(clknet_1_1__leaf__04623_),
    .D(net1428),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12063_ (.CLK(clknet_1_1__leaf__04623_),
    .D(net1421),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12064_ (.CLK(clknet_1_0__leaf__04623_),
    .D(net1289),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12065_ (.CLK(clknet_1_1__leaf__04623_),
    .D(net1646),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12066_ (.CLK(clknet_1_0__leaf__04623_),
    .D(net1639),
    .RESET_B(net823),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12067_ (.CLK(clknet_1_0__leaf__04623_),
    .D(net1631),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12068_ (.CLK(clknet_1_1__leaf__04623_),
    .D(net1624),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12069_ (.CLK(clknet_1_0__leaf__04623_),
    .D(net1617),
    .RESET_B(net823),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12070_ (.CLK(clknet_1_0__leaf__04622_),
    .D(net1295),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12071_ (.CLK(clknet_1_0__leaf__04622_),
    .D(net1573),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12072_ (.CLK(clknet_1_0__leaf__04622_),
    .D(net1492),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12073_ (.CLK(clknet_1_0__leaf__04622_),
    .D(net1468),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12074_ (.CLK(clknet_1_1__leaf__04622_),
    .D(net1459),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12075_ (.CLK(clknet_1_1__leaf__04622_),
    .D(net1451),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12076_ (.CLK(clknet_1_1__leaf__04622_),
    .D(net1443),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12077_ (.CLK(clknet_1_1__leaf__04622_),
    .D(net1435),
    .RESET_B(net840),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12078_ (.CLK(clknet_1_1__leaf__04621_),
    .D(net1536),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12079_ (.CLK(clknet_1_1__leaf__04621_),
    .D(net1528),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12080_ (.CLK(clknet_1_1__leaf__04621_),
    .D(net1521),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12081_ (.CLK(clknet_1_1__leaf__04621_),
    .D(net1514),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12082_ (.CLK(clknet_1_0__leaf__04621_),
    .D(net1507),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12083_ (.CLK(clknet_1_0__leaf__04621_),
    .D(net1502),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12084_ (.CLK(clknet_1_0__leaf__04621_),
    .D(net1483),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12085_ (.CLK(clknet_1_0__leaf__04621_),
    .D(net1476),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12086_ (.CLK(clknet_1_0__leaf__04620_),
    .D(net1605),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12087_ (.CLK(clknet_1_0__leaf__04620_),
    .D(net1597),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12088_ (.CLK(clknet_1_0__leaf__04620_),
    .D(net1594),
    .RESET_B(net819),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12089_ (.CLK(clknet_1_1__leaf__04620_),
    .D(net1580),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12090_ (.CLK(clknet_1_1__leaf__04620_),
    .D(net1565),
    .RESET_B(net830),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12091_ (.CLK(clknet_1_1__leaf__04620_),
    .D(net1558),
    .RESET_B(net830),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12092_ (.CLK(clknet_1_1__leaf__04620_),
    .D(net1551),
    .RESET_B(net830),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12093_ (.CLK(clknet_1_0__leaf__04620_),
    .D(net1544),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.u_reg.reg_2[23] ));
 sky130_fd_sc_hd__dfrtp_2 _12094_ (.CLK(clknet_1_1__leaf__04627_),
    .D(net1428),
    .RESET_B(net827),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[8] ));
 sky130_fd_sc_hd__dfrtp_2 _12095_ (.CLK(clknet_1_1__leaf__04627_),
    .D(net1421),
    .RESET_B(net827),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[9] ));
 sky130_fd_sc_hd__dfrtp_2 _12096_ (.CLK(clknet_1_1__leaf__04627_),
    .D(net1289),
    .RESET_B(net826),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[10] ));
 sky130_fd_sc_hd__dfrtp_2 _12097_ (.CLK(clknet_1_0__leaf__04627_),
    .D(net1646),
    .RESET_B(net828),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12098_ (.CLK(clknet_1_0__leaf__04627_),
    .D(net1639),
    .RESET_B(net823),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[12] ));
 sky130_fd_sc_hd__dfrtp_2 _12099_ (.CLK(clknet_1_0__leaf__04627_),
    .D(net1631),
    .RESET_B(net822),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[13] ));
 sky130_fd_sc_hd__dfrtp_4 _12100_ (.CLK(clknet_1_1__leaf__04627_),
    .D(net1624),
    .RESET_B(net827),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12101_ (.CLK(clknet_1_0__leaf__04627_),
    .D(net1617),
    .RESET_B(net824),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12102_ (.CLK(clknet_1_1__leaf__04626_),
    .D(net1295),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12103_ (.CLK(clknet_1_1__leaf__04626_),
    .D(net1573),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[1] ));
 sky130_fd_sc_hd__dfrtp_2 _12104_ (.CLK(clknet_1_1__leaf__04626_),
    .D(net1492),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12105_ (.CLK(clknet_1_0__leaf__04626_),
    .D(net1468),
    .RESET_B(net837),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[3] ));
 sky130_fd_sc_hd__dfrtp_2 _12106_ (.CLK(clknet_1_0__leaf__04626_),
    .D(net1459),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12107_ (.CLK(clknet_1_1__leaf__04626_),
    .D(net1451),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12108_ (.CLK(clknet_1_0__leaf__04626_),
    .D(net1443),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12109_ (.CLK(clknet_1_0__leaf__04626_),
    .D(net1435),
    .RESET_B(net839),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp2[7] ));
 sky130_fd_sc_hd__dfrtp_2 _12110_ (.CLK(clknet_1_0__leaf__04625_),
    .D(net1536),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12111_ (.CLK(clknet_1_0__leaf__04625_),
    .D(net1528),
    .RESET_B(net756),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12112_ (.CLK(clknet_1_0__leaf__04625_),
    .D(net1521),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[10] ));
 sky130_fd_sc_hd__dfrtp_2 _12113_ (.CLK(clknet_1_0__leaf__04625_),
    .D(net1514),
    .RESET_B(net757),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[11] ));
 sky130_fd_sc_hd__dfrtp_2 _12114_ (.CLK(clknet_1_1__leaf__04625_),
    .D(net1509),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12115_ (.CLK(clknet_1_1__leaf__04625_),
    .D(net1502),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12116_ (.CLK(clknet_1_1__leaf__04625_),
    .D(net1483),
    .RESET_B(net760),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12117_ (.CLK(clknet_1_1__leaf__04625_),
    .D(net1476),
    .RESET_B(net761),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12118_ (.CLK(clknet_1_0__leaf__04624_),
    .D(net1612),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[0] ));
 sky130_fd_sc_hd__dfrtp_2 _12119_ (.CLK(clknet_1_0__leaf__04624_),
    .D(net1597),
    .RESET_B(net820),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12120_ (.CLK(clknet_1_0__leaf__04624_),
    .D(net1594),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[2] ));
 sky130_fd_sc_hd__dfrtp_2 _12121_ (.CLK(clknet_1_1__leaf__04624_),
    .D(net1580),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[3] ));
 sky130_fd_sc_hd__dfrtp_2 _12122_ (.CLK(clknet_1_1__leaf__04624_),
    .D(net1565),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[4] ));
 sky130_fd_sc_hd__dfrtp_2 _12123_ (.CLK(clknet_1_1__leaf__04624_),
    .D(net111),
    .RESET_B(net831),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12124_ (.CLK(clknet_1_1__leaf__04624_),
    .D(net1551),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12125_ (.CLK(clknet_1_0__leaf__04624_),
    .D(net1544),
    .RESET_B(net829),
    .Q(\u_pwm.u_pwm_2.cfg_pwm_comp3[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12126_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[0] ),
    .RESET_B(net845),
    .Q(\u_pwm.reg_rdata_pwm2[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12127_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[1] ),
    .RESET_B(net845),
    .Q(\u_pwm.reg_rdata_pwm2[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12128_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[2] ),
    .RESET_B(net845),
    .Q(\u_pwm.reg_rdata_pwm2[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12129_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[3] ),
    .RESET_B(net846),
    .Q(\u_pwm.reg_rdata_pwm2[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12130_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[4] ),
    .RESET_B(net846),
    .Q(\u_pwm.reg_rdata_pwm2[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12131_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[5] ),
    .RESET_B(net845),
    .Q(\u_pwm.reg_rdata_pwm2[5] ));
 sky130_fd_sc_hd__dfrtp_2 _12132_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[6] ),
    .RESET_B(net844),
    .Q(\u_pwm.reg_rdata_pwm2[6] ));
 sky130_fd_sc_hd__dfrtp_2 _12133_ (.CLK(clknet_2_2__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[7] ),
    .RESET_B(net843),
    .Q(\u_pwm.reg_rdata_pwm2[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12134_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[8] ),
    .RESET_B(net834),
    .Q(\u_pwm.reg_rdata_pwm2[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12135_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[9] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12136_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[10] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12137_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[11] ),
    .RESET_B(net853),
    .Q(\u_pwm.reg_rdata_pwm2[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12138_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[12] ),
    .RESET_B(net853),
    .Q(\u_pwm.reg_rdata_pwm2[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12139_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[13] ),
    .RESET_B(net852),
    .Q(\u_pwm.reg_rdata_pwm2[13] ));
 sky130_fd_sc_hd__dfrtp_2 _12140_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[14] ),
    .RESET_B(net853),
    .Q(\u_pwm.reg_rdata_pwm2[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12141_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[15] ),
    .RESET_B(net827),
    .Q(\u_pwm.reg_rdata_pwm2[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12142_ (.CLK(clknet_2_3__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[16] ),
    .RESET_B(net831),
    .Q(\u_pwm.reg_rdata_pwm2[16] ));
 sky130_fd_sc_hd__dfrtp_1 _12143_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[17] ),
    .RESET_B(net834),
    .Q(\u_pwm.reg_rdata_pwm2[17] ));
 sky130_fd_sc_hd__dfrtp_1 _12144_ (.CLK(clknet_2_3__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[18] ),
    .RESET_B(net831),
    .Q(\u_pwm.reg_rdata_pwm2[18] ));
 sky130_fd_sc_hd__dfrtp_1 _12145_ (.CLK(clknet_2_3__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[19] ),
    .RESET_B(net831),
    .Q(\u_pwm.reg_rdata_pwm2[19] ));
 sky130_fd_sc_hd__dfrtp_1 _12146_ (.CLK(clknet_2_3__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[20] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[20] ));
 sky130_fd_sc_hd__dfrtp_1 _12147_ (.CLK(clknet_2_3__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[21] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[21] ));
 sky130_fd_sc_hd__dfrtp_1 _12148_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[22] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[22] ));
 sky130_fd_sc_hd__dfrtp_1 _12149_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[23] ),
    .RESET_B(net832),
    .Q(\u_pwm.reg_rdata_pwm2[23] ));
 sky130_fd_sc_hd__dfrtp_1 _12150_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[24] ),
    .RESET_B(net828),
    .Q(\u_pwm.reg_rdata_pwm2[24] ));
 sky130_fd_sc_hd__dfrtp_1 _12151_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[25] ),
    .RESET_B(net769),
    .Q(\u_pwm.reg_rdata_pwm2[25] ));
 sky130_fd_sc_hd__dfrtp_1 _12152_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[26] ),
    .RESET_B(net828),
    .Q(\u_pwm.reg_rdata_pwm2[26] ));
 sky130_fd_sc_hd__dfrtp_1 _12153_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[27] ),
    .RESET_B(net769),
    .Q(\u_pwm.reg_rdata_pwm2[27] ));
 sky130_fd_sc_hd__dfrtp_1 _12154_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[28] ),
    .RESET_B(net852),
    .Q(\u_pwm.reg_rdata_pwm2[28] ));
 sky130_fd_sc_hd__dfrtp_1 _12155_ (.CLK(clknet_2_0__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[29] ),
    .RESET_B(net767),
    .Q(\u_pwm.reg_rdata_pwm2[29] ));
 sky130_fd_sc_hd__dfrtp_1 _12156_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[30] ),
    .RESET_B(net828),
    .Q(\u_pwm.reg_rdata_pwm2[30] ));
 sky130_fd_sc_hd__dfrtp_1 _12157_ (.CLK(clknet_2_1__leaf__04608_),
    .D(\u_pwm.u_pwm_2.u_reg.reg_out[31] ),
    .RESET_B(net796),
    .Q(\u_pwm.reg_rdata_pwm2[31] ));
 sky130_fd_sc_hd__dfrtp_1 _12158_ (.CLK(clknet_4_12__leaf_mclk),
    .D(_00458_),
    .RESET_B(net977),
    .Q(\u_pwm.reg_ack_pwm2 ));
 sky130_fd_sc_hd__dfrtp_2 _12159_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00425_),
    .RESET_B(net821),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[0] ));
 sky130_fd_sc_hd__dfrtp_4 _12160_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00432_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[1] ));
 sky130_fd_sc_hd__dfrtp_4 _12161_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00433_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[2] ));
 sky130_fd_sc_hd__dfrtp_4 _12162_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00434_),
    .RESET_B(net821),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[3] ));
 sky130_fd_sc_hd__dfrtp_4 _12163_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00435_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[4] ));
 sky130_fd_sc_hd__dfrtp_4 _12164_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00436_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[5] ));
 sky130_fd_sc_hd__dfrtp_4 _12165_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00437_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[6] ));
 sky130_fd_sc_hd__dfrtp_4 _12166_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00438_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[7] ));
 sky130_fd_sc_hd__dfrtp_4 _12167_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00439_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[8] ));
 sky130_fd_sc_hd__dfrtp_4 _12168_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00440_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12169_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00426_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[10] ));
 sky130_fd_sc_hd__dfrtp_4 _12170_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00427_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[11] ));
 sky130_fd_sc_hd__dfrtp_4 _12171_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00428_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[12] ));
 sky130_fd_sc_hd__dfrtp_4 _12172_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00429_),
    .RESET_B(net816),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12173_ (.CLK(clknet_1_0__leaf__04606_),
    .D(_00430_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[14] ));
 sky130_fd_sc_hd__dfrtp_1 _12174_ (.CLK(clknet_1_1__leaf__04606_),
    .D(_00431_),
    .RESET_B(net818),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[15] ));
 sky130_fd_sc_hd__dfrtp_1 _12175_ (.CLK(_04607_),
    .D(\u_pwm.u_pwm_2.u_pwm.pwm_wfm_i ),
    .RESET_B(net852),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_wfm_r ));
 sky130_fd_sc_hd__dfrtp_1 _12176_ (.CLK(clknet_leaf_96_mclk),
    .D(\u_pwm.u_pwm_2.u_pwm.pwm_ovflow ),
    .RESET_B(net835),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_ovflow_l ));
 sky130_fd_sc_hd__dfrtp_1 _12177_ (.CLK(clknet_leaf_96_mclk),
    .D(_00424_),
    .RESET_B(net844),
    .Q(\u_pwm.u_pwm_2.gpio_tgr ));
 sky130_fd_sc_hd__dfrtp_1 _12178_ (.CLK(clknet_leaf_96_mclk),
    .D(_00423_),
    .RESET_B(net843),
    .Q(\u_pwm.u_pwm_2.u_pwm.gpio_l ));
 sky130_fd_sc_hd__dfrtp_1 _12179_ (.CLK(clknet_leaf_95_mclk),
    .D(_00441_),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[0] ));
 sky130_fd_sc_hd__dfrtp_1 _12180_ (.CLK(clknet_leaf_95_mclk),
    .D(_00447_),
    .RESET_B(net845),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[1] ));
 sky130_fd_sc_hd__dfrtp_1 _12181_ (.CLK(clknet_leaf_95_mclk),
    .D(_00448_),
    .RESET_B(net851),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[2] ));
 sky130_fd_sc_hd__dfrtp_1 _12182_ (.CLK(clknet_leaf_95_mclk),
    .D(_00449_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[3] ));
 sky130_fd_sc_hd__dfrtp_1 _12183_ (.CLK(clknet_leaf_93_mclk),
    .D(_00450_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[4] ));
 sky130_fd_sc_hd__dfrtp_1 _12184_ (.CLK(clknet_leaf_93_mclk),
    .D(_00451_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[5] ));
 sky130_fd_sc_hd__dfrtp_1 _12185_ (.CLK(clknet_leaf_93_mclk),
    .D(_00452_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[6] ));
 sky130_fd_sc_hd__dfrtp_1 _12186_ (.CLK(clknet_leaf_93_mclk),
    .D(_00453_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[7] ));
 sky130_fd_sc_hd__dfrtp_1 _12187_ (.CLK(clknet_leaf_93_mclk),
    .D(_00454_),
    .RESET_B(net841),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[8] ));
 sky130_fd_sc_hd__dfrtp_1 _12188_ (.CLK(clknet_leaf_93_mclk),
    .D(_00455_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[9] ));
 sky130_fd_sc_hd__dfrtp_1 _12189_ (.CLK(clknet_leaf_94_mclk),
    .D(_00442_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[10] ));
 sky130_fd_sc_hd__dfrtp_1 _12190_ (.CLK(clknet_leaf_93_mclk),
    .D(_00443_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[11] ));
 sky130_fd_sc_hd__dfrtp_1 _12191_ (.CLK(clknet_leaf_93_mclk),
    .D(_00444_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[12] ));
 sky130_fd_sc_hd__dfrtp_1 _12192_ (.CLK(clknet_leaf_93_mclk),
    .D(_00445_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[13] ));
 sky130_fd_sc_hd__dfrtp_1 _12193_ (.CLK(clknet_leaf_93_mclk),
    .D(_00446_),
    .RESET_B(net838),
    .Q(\u_pwm.u_pwm_2.u_pwm.pwm_scnt[14] ));
 sky130_fd_sc_hd__clkbuf_1 _12231_ (.A(\u_glbl_reg.reg_2[16] ),
    .X(net232));
 sky130_fd_sc_hd__clkbuf_1 _12232_ (.A(\u_glbl_reg.reg_2[17] ),
    .X(net239));
 sky130_fd_sc_hd__clkbuf_1 _12233_ (.A(\u_glbl_reg.reg_2[18] ),
    .X(net240));
 sky130_fd_sc_hd__clkbuf_1 _12234_ (.A(\u_glbl_reg.reg_2[19] ),
    .X(net241));
 sky130_fd_sc_hd__clkbuf_1 _12235_ (.A(\u_glbl_reg.reg_2[20] ),
    .X(net242));
 sky130_fd_sc_hd__clkbuf_1 _12236_ (.A(\u_glbl_reg.reg_2[21] ),
    .X(net243));
 sky130_fd_sc_hd__clkbuf_1 _12237_ (.A(\u_glbl_reg.reg_2[22] ),
    .X(net244));
 sky130_fd_sc_hd__clkbuf_1 _12238_ (.A(\u_glbl_reg.reg_2[23] ),
    .X(net245));
 sky130_fd_sc_hd__clkbuf_1 _12239_ (.A(\u_glbl_reg.reg_2[24] ),
    .X(net246));
 sky130_fd_sc_hd__clkbuf_1 _12240_ (.A(\u_glbl_reg.reg_2[25] ),
    .X(net247));
 sky130_fd_sc_hd__clkbuf_1 _12241_ (.A(\u_glbl_reg.reg_2[26] ),
    .X(net233));
 sky130_fd_sc_hd__clkbuf_1 _12242_ (.A(\u_glbl_reg.reg_2[27] ),
    .X(net234));
 sky130_fd_sc_hd__clkbuf_1 _12243_ (.A(\u_glbl_reg.reg_2[28] ),
    .X(net235));
 sky130_fd_sc_hd__clkbuf_1 _12244_ (.A(\u_glbl_reg.reg_2[29] ),
    .X(net236));
 sky130_fd_sc_hd__clkbuf_1 _12245_ (.A(\u_glbl_reg.reg_2[30] ),
    .X(net237));
 sky130_fd_sc_hd__clkbuf_1 _12246_ (.A(\u_glbl_reg.reg_2[31] ),
    .X(net238));
 sky130_fd_sc_hd__clkbuf_1 _12247_ (.A(\u_glbl_reg.u_buf_cpu0_rst.X ),
    .X(net248));
 sky130_fd_sc_hd__clkbuf_1 _12248_ (.A(\u_glbl_reg.u_buf_cpu1_rst.X ),
    .X(net249));
 sky130_fd_sc_hd__clkbuf_1 _12249_ (.A(\u_glbl_reg.u_buf_cpu2_rst.X ),
    .X(net250));
 sky130_fd_sc_hd__clkbuf_1 _12250_ (.A(\u_glbl_reg.u_buf_cpu3_rst.X ),
    .X(net251));
 sky130_fd_sc_hd__clkbuf_1 _12251_ (.A(net1652),
    .X(net273));
 sky130_fd_sc_hd__clkbuf_1 _12252_ (.A(net1652),
    .X(net274));
 sky130_fd_sc_hd__clkbuf_1 _12253_ (.A(net1652),
    .X(net276));
 sky130_fd_sc_hd__clkbuf_1 _12254_ (.A(net1652),
    .X(net277));
 sky130_fd_sc_hd__clkbuf_1 _12255_ (.A(net1653),
    .X(net278));
 sky130_fd_sc_hd__clkbuf_1 _12256_ (.A(net1653),
    .X(net283));
 sky130_fd_sc_hd__buf_4 _12257_ (.A(net143),
    .X(net311));
 sky130_fd_sc_hd__buf_4 _12258_ (.A(net144),
    .X(net312));
 sky130_fd_sc_hd__buf_4 _12259_ (.A(net145),
    .X(net314));
 sky130_fd_sc_hd__buf_4 _12260_ (.A(net146),
    .X(net315));
 sky130_fd_sc_hd__buf_4 _12261_ (.A(net147),
    .X(net316));
 sky130_fd_sc_hd__buf_4 _12262_ (.A(net135),
    .X(net317));
 sky130_fd_sc_hd__buf_4 _12263_ (.A(net136),
    .X(net318));
 sky130_fd_sc_hd__buf_4 _12264_ (.A(net137),
    .X(net319));
 sky130_fd_sc_hd__buf_4 _12265_ (.A(net138),
    .X(net320));
 sky130_fd_sc_hd__clkbuf_1 _12266_ (.A(\u_glbl_reg.dbg_clk_mon ),
    .X(net321));
 sky130_fd_sc_hd__clkbuf_1 _12267_ (.A(net1339),
    .X(net332));
 sky130_fd_sc_hd__clkbuf_2 _12268_ (.A(net1376),
    .X(net369));
 sky130_fd_sc_hd__clkbuf_2 _12269_ (.A(net1373),
    .X(net371));
 sky130_fd_sc_hd__clkbuf_1 _12270_ (.A(net1371),
    .X(net372));
 sky130_fd_sc_hd__clkbuf_2 _12271_ (.A(net1357),
    .X(net373));
 sky130_fd_sc_hd__clkbuf_2 _12272_ (.A(net1347),
    .X(net374));
 sky130_fd_sc_hd__clkbuf_2 _12273_ (.A(net1345),
    .X(net375));
 sky130_fd_sc_hd__clkbuf_2 _12274_ (.A(net1344),
    .X(net376));
 sky130_fd_sc_hd__clkbuf_1 _12275_ (.A(net1342),
    .X(net377));
 sky130_fd_sc_hd__clkbuf_1 _12276_ (.A(net1341),
    .X(net378));
 sky130_fd_sc_hd__clkbuf_1 _12277_ (.A(net1340),
    .X(net379));
 sky130_fd_sc_hd__clkbuf_1 _12278_ (.A(net1374),
    .X(net370));
 sky130_fd_sc_hd__clkbuf_1 _12279_ (.A(net1337),
    .X(net380));
 sky130_fd_sc_hd__clkbuf_1 _12280_ (.A(net1330),
    .X(net381));
 sky130_fd_sc_hd__clkbuf_1 _12281_ (.A(net1322),
    .X(net382));
 sky130_fd_sc_hd__clkbuf_1 _12282_ (.A(net1315),
    .X(net383));
 sky130_fd_sc_hd__clkbuf_1 _12283_ (.A(net1302),
    .X(net385));
 sky130_fd_sc_hd__clkbuf_1 _12284_ (.A(net1576),
    .X(net396));
 sky130_fd_sc_hd__clkbuf_1 _12285_ (.A(net1495),
    .X(net407));
 sky130_fd_sc_hd__clkbuf_1 _12286_ (.A(net1472),
    .X(net410));
 sky130_fd_sc_hd__clkbuf_1 _12287_ (.A(net1462),
    .X(net411));
 sky130_fd_sc_hd__clkbuf_1 _12288_ (.A(net1454),
    .X(net412));
 sky130_fd_sc_hd__clkbuf_1 _12289_ (.A(net1446),
    .X(net413));
 sky130_fd_sc_hd__clkbuf_1 _12290_ (.A(net1437),
    .X(net414));
 sky130_fd_sc_hd__clkbuf_1 _12291_ (.A(net1431),
    .X(net415));
 sky130_fd_sc_hd__clkbuf_1 _12292_ (.A(net1424),
    .X(net416));
 sky130_fd_sc_hd__clkbuf_1 _12293_ (.A(net1292),
    .X(net386));
 sky130_fd_sc_hd__clkbuf_1 _12294_ (.A(net1649),
    .X(net387));
 sky130_fd_sc_hd__clkbuf_1 _12295_ (.A(net1642),
    .X(net388));
 sky130_fd_sc_hd__clkbuf_1 _12296_ (.A(net1634),
    .X(net389));
 sky130_fd_sc_hd__clkbuf_1 _12297_ (.A(net1627),
    .X(net390));
 sky130_fd_sc_hd__clkbuf_1 _12298_ (.A(net1620),
    .X(net391));
 sky130_fd_sc_hd__clkbuf_1 _12299_ (.A(net1609),
    .X(net392));
 sky130_fd_sc_hd__clkbuf_1 _12300_ (.A(net1601),
    .X(net393));
 sky130_fd_sc_hd__clkbuf_1 _12301_ (.A(net1593),
    .X(net394));
 sky130_fd_sc_hd__clkbuf_1 _12302_ (.A(net1585),
    .X(net395));
 sky130_fd_sc_hd__clkbuf_1 _12303_ (.A(net1570),
    .X(net397));
 sky130_fd_sc_hd__clkbuf_1 _12304_ (.A(net1563),
    .X(net398));
 sky130_fd_sc_hd__clkbuf_1 _12305_ (.A(net1554),
    .X(net399));
 sky130_fd_sc_hd__clkbuf_1 _12306_ (.A(net1548),
    .X(net400));
 sky130_fd_sc_hd__clkbuf_1 _12307_ (.A(net1540),
    .X(net401));
 sky130_fd_sc_hd__clkbuf_1 _12308_ (.A(net1532),
    .X(net402));
 sky130_fd_sc_hd__clkbuf_1 _12309_ (.A(net1525),
    .X(net403));
 sky130_fd_sc_hd__clkbuf_1 _12310_ (.A(net1518),
    .X(net404));
 sky130_fd_sc_hd__clkbuf_1 _12311_ (.A(net1511),
    .X(net405));
 sky130_fd_sc_hd__clkbuf_1 _12312_ (.A(net1504),
    .X(net406));
 sky130_fd_sc_hd__clkbuf_1 _12313_ (.A(net1487),
    .X(net408));
 sky130_fd_sc_hd__clkbuf_1 _12314_ (.A(net1480),
    .X(net409));
 sky130_fd_sc_hd__clkbuf_1 _12315_ (.A(net1416),
    .X(net417));
 sky130_fd_sc_hd__clkbuf_1 _12316_ (.A(net1395),
    .X(net455));
 sky130_fd_sc_hd__clkbuf_1 _12317_ (.A(net1393),
    .X(net456));
 sky130_fd_sc_hd__clkbuf_4 _12318_ (.A(net1391),
    .X(net457));
 sky130_fd_sc_hd__clkbuf_1 _12319_ (.A(net1389),
    .X(net458));
 sky130_fd_sc_hd__clkbuf_1 _12320_ (.A(\u_glbl_reg.reg_12[13] ),
    .X(net497));
 sky130_fd_sc_hd__clkbuf_1 _12321_ (.A(\u_glbl_reg.reg_12[14] ),
    .X(net498));
 sky130_fd_sc_hd__clkbuf_1 _12322_ (.A(\u_glbl_reg.u_buf_uart0_rst.X ),
    .X(net499));
 sky130_fd_sc_hd__clkbuf_1 _12323_ (.A(\u_glbl_reg.u_buf_uart1_rst.X ),
    .X(net500));
 sky130_fd_sc_hd__clkbuf_1 _12324_ (.A(\u_glbl_reg.reg_2[0] ),
    .X(net508));
 sky130_fd_sc_hd__clkbuf_2 _12325_ (.A(\u_glbl_reg.reg_2[1] ),
    .X(net509));
 sky130_fd_sc_hd__clkbuf_1 _12326_ (.A(\u_glbl_reg.reg_2[2] ),
    .X(net510));
 sky130_fd_sc_hd__clkbuf_1 _12327_ (.A(net1375),
    .X(net512));
 sky130_fd_sc_hd__dlclkp_4 _12328_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00038_),
    .GCLK(_04353_));
 sky130_fd_sc_hd__dlclkp_1 _12329_ (.CLK(\u_glbl_reg.dbg_clk_ref_buf ),
    .GATE(_00044_),
    .GCLK(_04354_));
 sky130_fd_sc_hd__dlclkp_1 _12330_ (.CLK(\u_glbl_reg.dbg_clk_ref_buf ),
    .GATE(_00045_),
    .GCLK(_04355_));
 sky130_fd_sc_hd__dlclkp_1 _12331_ (.CLK(clknet_1_1__leaf_user_clock1),
    .GATE(_00054_),
    .GCLK(_04356_));
 sky130_fd_sc_hd__dlclkp_1 _12332_ (.CLK(clknet_1_1__leaf_user_clock1),
    .GATE(_00055_),
    .GCLK(_04357_));
 sky130_fd_sc_hd__dlclkp_4 _12333_ (.CLK(clknet_leaf_33_mclk),
    .GATE(\u_glbl_reg.reg_ack ),
    .GCLK(_04358_));
 sky130_fd_sc_hd__dlclkp_4 _12334_ (.CLK(clknet_leaf_33_mclk),
    .GATE(\u_glbl_reg.reg_ack ),
    .GCLK(_04359_));
 sky130_fd_sc_hd__dlclkp_1 _12335_ (.CLK(clknet_leaf_19_mclk),
    .GATE(_00059_),
    .GCLK(_04360_));
 sky130_fd_sc_hd__dlclkp_1 _12336_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00060_),
    .GCLK(_04361_));
 sky130_fd_sc_hd__dlclkp_1 _12337_ (.CLK(clknet_leaf_13_mclk),
    .GATE(_00061_),
    .GCLK(_04362_));
 sky130_fd_sc_hd__dlclkp_1 _12338_ (.CLK(clknet_leaf_9_mclk),
    .GATE(_00062_),
    .GCLK(_04363_));
 sky130_fd_sc_hd__dlclkp_1 _12339_ (.CLK(clknet_leaf_9_mclk),
    .GATE(_00063_),
    .GCLK(_04364_));
 sky130_fd_sc_hd__dlclkp_1 _12340_ (.CLK(clknet_leaf_9_mclk),
    .GATE(_00064_),
    .GCLK(_04365_));
 sky130_fd_sc_hd__dlclkp_1 _12341_ (.CLK(clknet_leaf_8_mclk),
    .GATE(_00065_),
    .GCLK(_04366_));
 sky130_fd_sc_hd__dlclkp_1 _12342_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00066_),
    .GCLK(_04367_));
 sky130_fd_sc_hd__dlclkp_1 _12343_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00067_),
    .GCLK(_04368_));
 sky130_fd_sc_hd__dlclkp_1 _12344_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00068_),
    .GCLK(_04369_));
 sky130_fd_sc_hd__dlclkp_1 _12345_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00069_),
    .GCLK(_04370_));
 sky130_fd_sc_hd__dlclkp_1 _12346_ (.CLK(clknet_leaf_25_mclk),
    .GATE(_00070_),
    .GCLK(_04371_));
 sky130_fd_sc_hd__dlclkp_1 _12347_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00071_),
    .GCLK(_04372_));
 sky130_fd_sc_hd__dlclkp_1 _12348_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00072_),
    .GCLK(_04373_));
 sky130_fd_sc_hd__dlclkp_1 _12349_ (.CLK(clknet_leaf_26_mclk),
    .GATE(_00073_),
    .GCLK(_04374_));
 sky130_fd_sc_hd__dlclkp_1 _12350_ (.CLK(clknet_leaf_24_mclk),
    .GATE(_00074_),
    .GCLK(_04375_));
 sky130_fd_sc_hd__dlclkp_1 _12351_ (.CLK(clknet_leaf_110_mclk),
    .GATE(_00075_),
    .GCLK(_04376_));
 sky130_fd_sc_hd__dlclkp_1 _12352_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00076_),
    .GCLK(_04377_));
 sky130_fd_sc_hd__dlclkp_1 _12353_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00077_),
    .GCLK(_04378_));
 sky130_fd_sc_hd__dlclkp_1 _12354_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00078_),
    .GCLK(_04379_));
 sky130_fd_sc_hd__dlclkp_1 _12355_ (.CLK(clknet_leaf_110_mclk),
    .GATE(_00079_),
    .GCLK(_04380_));
 sky130_fd_sc_hd__dlclkp_1 _12356_ (.CLK(clknet_leaf_110_mclk),
    .GATE(_00080_),
    .GCLK(_04381_));
 sky130_fd_sc_hd__dlclkp_1 _12357_ (.CLK(clknet_leaf_19_mclk),
    .GATE(_00081_),
    .GCLK(_04382_));
 sky130_fd_sc_hd__dlclkp_1 _12358_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00082_),
    .GCLK(_04383_));
 sky130_fd_sc_hd__dlclkp_1 _12359_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00083_),
    .GCLK(_04384_));
 sky130_fd_sc_hd__dlclkp_1 _12360_ (.CLK(clknet_leaf_10_mclk),
    .GATE(_00084_),
    .GCLK(_04385_));
 sky130_fd_sc_hd__dlclkp_1 _12361_ (.CLK(clknet_leaf_10_mclk),
    .GATE(_00085_),
    .GCLK(_04386_));
 sky130_fd_sc_hd__dlclkp_1 _12362_ (.CLK(clknet_leaf_13_mclk),
    .GATE(_00086_),
    .GCLK(_04387_));
 sky130_fd_sc_hd__dlclkp_1 _12363_ (.CLK(clknet_leaf_25_mclk),
    .GATE(_00087_),
    .GCLK(_04388_));
 sky130_fd_sc_hd__dlclkp_1 _12364_ (.CLK(clknet_leaf_25_mclk),
    .GATE(_00088_),
    .GCLK(_04389_));
 sky130_fd_sc_hd__dlclkp_1 _12365_ (.CLK(clknet_leaf_8_mclk),
    .GATE(_00089_),
    .GCLK(_04390_));
 sky130_fd_sc_hd__dlclkp_1 _12366_ (.CLK(clknet_leaf_9_mclk),
    .GATE(_00090_),
    .GCLK(_04391_));
 sky130_fd_sc_hd__dlclkp_2 _12367_ (.CLK(clknet_leaf_126_mclk),
    .GATE(_00123_),
    .GCLK(_04392_));
 sky130_fd_sc_hd__dlclkp_2 _12368_ (.CLK(clknet_leaf_7_mclk),
    .GATE(_00124_),
    .GCLK(_04393_));
 sky130_fd_sc_hd__dlclkp_2 _12369_ (.CLK(clknet_leaf_6_mclk),
    .GATE(_00125_),
    .GCLK(_04394_));
 sky130_fd_sc_hd__dlclkp_2 _12370_ (.CLK(clknet_leaf_126_mclk),
    .GATE(_00126_),
    .GCLK(_04395_));
 sky130_fd_sc_hd__dlclkp_2 _12371_ (.CLK(clknet_leaf_29_mclk),
    .GATE(_00127_),
    .GCLK(_04396_));
 sky130_fd_sc_hd__dlclkp_2 _12372_ (.CLK(clknet_leaf_128_mclk),
    .GATE(_00128_),
    .GCLK(_04397_));
 sky130_fd_sc_hd__dlclkp_2 _12373_ (.CLK(clknet_leaf_124_mclk),
    .GATE(_00129_),
    .GCLK(_04398_));
 sky130_fd_sc_hd__dlclkp_2 _12374_ (.CLK(clknet_leaf_5_mclk),
    .GATE(_00130_),
    .GCLK(_04399_));
 sky130_fd_sc_hd__dlclkp_2 _12375_ (.CLK(clknet_4_1__leaf_mclk),
    .GATE(_00131_),
    .GCLK(_04400_));
 sky130_fd_sc_hd__dlclkp_2 _12376_ (.CLK(clknet_leaf_25_mclk),
    .GATE(_00132_),
    .GCLK(_04401_));
 sky130_fd_sc_hd__dlclkp_2 _12377_ (.CLK(clknet_leaf_28_mclk),
    .GATE(_00133_),
    .GCLK(_04402_));
 sky130_fd_sc_hd__dlclkp_2 _12378_ (.CLK(clknet_leaf_4_mclk),
    .GATE(_00134_),
    .GCLK(_04403_));
 sky130_fd_sc_hd__dlclkp_2 _12379_ (.CLK(clknet_leaf_28_mclk),
    .GATE(_00135_),
    .GCLK(_04404_));
 sky130_fd_sc_hd__dlclkp_2 _12380_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00136_),
    .GCLK(_04405_));
 sky130_fd_sc_hd__dlclkp_2 _12381_ (.CLK(clknet_4_8__leaf_mclk),
    .GATE(_00137_),
    .GCLK(_04406_));
 sky130_fd_sc_hd__dlclkp_2 _12382_ (.CLK(clknet_leaf_122_mclk),
    .GATE(_00138_),
    .GCLK(_04407_));
 sky130_fd_sc_hd__dlclkp_2 _12383_ (.CLK(clknet_leaf_26_mclk),
    .GATE(_00139_),
    .GCLK(_04408_));
 sky130_fd_sc_hd__dlclkp_2 _12384_ (.CLK(clknet_leaf_126_mclk),
    .GATE(_00140_),
    .GCLK(_04409_));
 sky130_fd_sc_hd__dlclkp_2 _12385_ (.CLK(clknet_leaf_6_mclk),
    .GATE(_00141_),
    .GCLK(_04410_));
 sky130_fd_sc_hd__dlclkp_2 _12386_ (.CLK(clknet_leaf_122_mclk),
    .GATE(_00142_),
    .GCLK(_04411_));
 sky130_fd_sc_hd__dlclkp_2 _12387_ (.CLK(clknet_leaf_31_mclk),
    .GATE(_00143_),
    .GCLK(_04412_));
 sky130_fd_sc_hd__dlclkp_2 _12388_ (.CLK(clknet_leaf_2_mclk),
    .GATE(_00144_),
    .GCLK(_04413_));
 sky130_fd_sc_hd__dlclkp_2 _12389_ (.CLK(clknet_leaf_123_mclk),
    .GATE(_00145_),
    .GCLK(_04414_));
 sky130_fd_sc_hd__dlclkp_2 _12390_ (.CLK(clknet_leaf_7_mclk),
    .GATE(_00146_),
    .GCLK(_04415_));
 sky130_fd_sc_hd__dlclkp_2 _12391_ (.CLK(clknet_leaf_124_mclk),
    .GATE(_00147_),
    .GCLK(_04416_));
 sky130_fd_sc_hd__dlclkp_2 _12392_ (.CLK(clknet_leaf_5_mclk),
    .GATE(_00148_),
    .GCLK(_04417_));
 sky130_fd_sc_hd__dlclkp_2 _12393_ (.CLK(clknet_leaf_4_mclk),
    .GATE(_00149_),
    .GCLK(_04418_));
 sky130_fd_sc_hd__dlclkp_2 _12394_ (.CLK(clknet_leaf_128_mclk),
    .GATE(_00150_),
    .GCLK(_04419_));
 sky130_fd_sc_hd__dlclkp_2 _12395_ (.CLK(clknet_leaf_29_mclk),
    .GATE(_00151_),
    .GCLK(_04420_));
 sky130_fd_sc_hd__dlclkp_2 _12396_ (.CLK(clknet_leaf_123_mclk),
    .GATE(_00152_),
    .GCLK(_04421_));
 sky130_fd_sc_hd__dlclkp_2 _12397_ (.CLK(clknet_leaf_120_mclk),
    .GATE(_00153_),
    .GCLK(_04422_));
 sky130_fd_sc_hd__dlclkp_2 _12398_ (.CLK(clknet_leaf_8_mclk),
    .GATE(_00154_),
    .GCLK(_04423_));
 sky130_fd_sc_hd__dlclkp_2 _12399_ (.CLK(clknet_leaf_29_mclk),
    .GATE(_00155_),
    .GCLK(_04424_));
 sky130_fd_sc_hd__dlclkp_2 _12400_ (.CLK(clknet_leaf_126_mclk),
    .GATE(_00156_),
    .GCLK(_04425_));
 sky130_fd_sc_hd__dlclkp_2 _12401_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00157_),
    .GCLK(_04426_));
 sky130_fd_sc_hd__dlclkp_2 _12402_ (.CLK(clknet_leaf_8_mclk),
    .GATE(_00158_),
    .GCLK(_04427_));
 sky130_fd_sc_hd__dlclkp_2 _12403_ (.CLK(clknet_leaf_30_mclk),
    .GATE(_00159_),
    .GCLK(_04428_));
 sky130_fd_sc_hd__dlclkp_2 _12404_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00160_),
    .GCLK(_04429_));
 sky130_fd_sc_hd__dlclkp_2 _12405_ (.CLK(clknet_leaf_122_mclk),
    .GATE(_00161_),
    .GCLK(_04430_));
 sky130_fd_sc_hd__dlclkp_2 _12406_ (.CLK(clknet_leaf_7_mclk),
    .GATE(_00162_),
    .GCLK(_04431_));
 sky130_fd_sc_hd__dlclkp_2 _12407_ (.CLK(clknet_leaf_6_mclk),
    .GATE(_00163_),
    .GCLK(_04432_));
 sky130_fd_sc_hd__dlclkp_2 _12408_ (.CLK(clknet_leaf_128_mclk),
    .GATE(_00164_),
    .GCLK(_04433_));
 sky130_fd_sc_hd__dlclkp_2 _12409_ (.CLK(clknet_leaf_124_mclk),
    .GATE(_00165_),
    .GCLK(_04434_));
 sky130_fd_sc_hd__dlclkp_2 _12410_ (.CLK(clknet_leaf_5_mclk),
    .GATE(_00166_),
    .GCLK(_04435_));
 sky130_fd_sc_hd__dlclkp_2 _12411_ (.CLK(clknet_leaf_28_mclk),
    .GATE(_00167_),
    .GCLK(_04436_));
 sky130_fd_sc_hd__dlclkp_2 _12412_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00168_),
    .GCLK(_04437_));
 sky130_fd_sc_hd__dlclkp_2 _12413_ (.CLK(clknet_leaf_10_mclk),
    .GATE(_00169_),
    .GCLK(_04438_));
 sky130_fd_sc_hd__dlclkp_2 _12414_ (.CLK(clknet_4_2__leaf_mclk),
    .GATE(_00170_),
    .GCLK(_04439_));
 sky130_fd_sc_hd__dlclkp_2 _12415_ (.CLK(clknet_leaf_112_mclk),
    .GATE(_00171_),
    .GCLK(_04440_));
 sky130_fd_sc_hd__dlclkp_2 _12416_ (.CLK(clknet_leaf_10_mclk),
    .GATE(_00172_),
    .GCLK(_04441_));
 sky130_fd_sc_hd__dlclkp_2 _12417_ (.CLK(clknet_leaf_26_mclk),
    .GATE(_00173_),
    .GCLK(_04442_));
 sky130_fd_sc_hd__dlclkp_2 _12418_ (.CLK(clknet_leaf_126_mclk),
    .GATE(_00174_),
    .GCLK(_04443_));
 sky130_fd_sc_hd__dlclkp_2 _12419_ (.CLK(clknet_leaf_5_mclk),
    .GATE(_00175_),
    .GCLK(_04444_));
 sky130_fd_sc_hd__dlclkp_2 _12420_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00176_),
    .GCLK(_04445_));
 sky130_fd_sc_hd__dlclkp_2 _12421_ (.CLK(clknet_4_0__leaf_mclk),
    .GATE(_00177_),
    .GCLK(_04446_));
 sky130_fd_sc_hd__dlclkp_2 _12422_ (.CLK(clknet_leaf_2_mclk),
    .GATE(_00178_),
    .GCLK(_04447_));
 sky130_fd_sc_hd__dlclkp_2 _12423_ (.CLK(clknet_leaf_7_mclk),
    .GATE(_00179_),
    .GCLK(_04448_));
 sky130_fd_sc_hd__dlclkp_2 _12424_ (.CLK(clknet_leaf_6_mclk),
    .GATE(_00180_),
    .GCLK(_04449_));
 sky130_fd_sc_hd__dlclkp_2 _12425_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00181_),
    .GCLK(_04450_));
 sky130_fd_sc_hd__dlclkp_2 _12426_ (.CLK(clknet_leaf_122_mclk),
    .GATE(_00182_),
    .GCLK(_04451_));
 sky130_fd_sc_hd__dlclkp_2 _12427_ (.CLK(clknet_leaf_47_mclk),
    .GATE(_00183_),
    .GCLK(_04452_));
 sky130_fd_sc_hd__dlclkp_2 _12428_ (.CLK(clknet_leaf_41_mclk),
    .GATE(_00184_),
    .GCLK(_04453_));
 sky130_fd_sc_hd__dlclkp_2 _12429_ (.CLK(clknet_leaf_43_mclk),
    .GATE(_00185_),
    .GCLK(_04454_));
 sky130_fd_sc_hd__dlclkp_2 _12430_ (.CLK(clknet_leaf_41_mclk),
    .GATE(_00186_),
    .GCLK(_04455_));
 sky130_fd_sc_hd__dlclkp_2 _12431_ (.CLK(\u_glbl_reg.rtc_ref_clk ),
    .GATE(_00193_),
    .GCLK(_04456_));
 sky130_fd_sc_hd__dlclkp_2 _12432_ (.CLK(\u_glbl_reg.rtc_ref_clk ),
    .GATE(_00194_),
    .GCLK(_04457_));
 sky130_fd_sc_hd__dlclkp_2 _12433_ (.CLK(clknet_leaf_122_mclk),
    .GATE(_00232_),
    .GCLK(_04458_));
 sky130_fd_sc_hd__dlclkp_2 _12434_ (.CLK(clknet_leaf_4_mclk),
    .GATE(_00233_),
    .GCLK(_04459_));
 sky130_fd_sc_hd__dlclkp_2 _12435_ (.CLK(clknet_leaf_1_mclk),
    .GATE(_00234_),
    .GCLK(_04460_));
 sky130_fd_sc_hd__dlclkp_2 _12436_ (.CLK(clknet_leaf_0_mclk),
    .GATE(_00235_),
    .GCLK(_04461_));
 sky130_fd_sc_hd__dlclkp_1 _12437_ (.CLK(clknet_leaf_0_mclk),
    .GATE(_00236_),
    .GCLK(_04462_));
 sky130_fd_sc_hd__dlclkp_2 _12438_ (.CLK(\u_glbl_reg.u_usb_clk_sel.A0 ),
    .GATE(_00243_),
    .GCLK(_04463_));
 sky130_fd_sc_hd__dlclkp_2 _12439_ (.CLK(\u_glbl_reg.u_usb_clk_sel.A0 ),
    .GATE(_00244_),
    .GCLK(_04464_));
 sky130_fd_sc_hd__dlclkp_1 _12440_ (.CLK(clknet_leaf_88_mclk),
    .GATE(_00250_),
    .GCLK(_04465_));
 sky130_fd_sc_hd__dlclkp_1 _12441_ (.CLK(clknet_leaf_110_mclk),
    .GATE(net720),
    .GCLK(_04466_));
 sky130_fd_sc_hd__dlclkp_1 _12442_ (.CLK(clknet_leaf_10_mclk),
    .GATE(net719),
    .GCLK(_04467_));
 sky130_fd_sc_hd__dlclkp_1 _12443_ (.CLK(clknet_leaf_15_mclk),
    .GATE(net719),
    .GCLK(_04468_));
 sky130_fd_sc_hd__dlclkp_1 _12444_ (.CLK(clknet_leaf_13_mclk),
    .GATE(net719),
    .GCLK(_04469_));
 sky130_fd_sc_hd__dlclkp_1 _12445_ (.CLK(clknet_leaf_8_mclk),
    .GATE(net722),
    .GCLK(_04470_));
 sky130_fd_sc_hd__dlclkp_1 _12446_ (.CLK(clknet_leaf_19_mclk),
    .GATE(net722),
    .GCLK(_04471_));
 sky130_fd_sc_hd__dlclkp_1 _12447_ (.CLK(clknet_leaf_75_mclk),
    .GATE(net722),
    .GCLK(_04472_));
 sky130_fd_sc_hd__dlclkp_1 _12448_ (.CLK(clknet_leaf_75_mclk),
    .GATE(net722),
    .GCLK(_04473_));
 sky130_fd_sc_hd__dlclkp_1 _12449_ (.CLK(clknet_leaf_24_mclk),
    .GATE(net722),
    .GCLK(_04474_));
 sky130_fd_sc_hd__dlclkp_1 _12450_ (.CLK(clknet_leaf_23_mclk),
    .GATE(net722),
    .GCLK(_04475_));
 sky130_fd_sc_hd__dlclkp_1 _12451_ (.CLK(clknet_leaf_107_mclk),
    .GATE(net719),
    .GCLK(_04476_));
 sky130_fd_sc_hd__dlclkp_1 _12452_ (.CLK(clknet_leaf_23_mclk),
    .GATE(net722),
    .GCLK(_04477_));
 sky130_fd_sc_hd__dlclkp_1 _12453_ (.CLK(clknet_leaf_23_mclk),
    .GATE(net722),
    .GCLK(_04478_));
 sky130_fd_sc_hd__dlclkp_1 _12454_ (.CLK(clknet_leaf_56_mclk),
    .GATE(net722),
    .GCLK(_04479_));
 sky130_fd_sc_hd__dlclkp_1 _12455_ (.CLK(clknet_leaf_115_mclk),
    .GATE(net719),
    .GCLK(_04480_));
 sky130_fd_sc_hd__dlclkp_1 _12456_ (.CLK(clknet_leaf_92_mclk),
    .GATE(net721),
    .GCLK(_04481_));
 sky130_fd_sc_hd__dlclkp_1 _12457_ (.CLK(clknet_leaf_114_mclk),
    .GATE(net719),
    .GCLK(_04482_));
 sky130_fd_sc_hd__dlclkp_1 _12458_ (.CLK(clknet_leaf_92_mclk),
    .GATE(net721),
    .GCLK(_04483_));
 sky130_fd_sc_hd__dlclkp_1 _12459_ (.CLK(clknet_leaf_91_mclk),
    .GATE(net721),
    .GCLK(_04484_));
 sky130_fd_sc_hd__dlclkp_1 _12460_ (.CLK(clknet_leaf_120_mclk),
    .GATE(net719),
    .GCLK(_04485_));
 sky130_fd_sc_hd__dlclkp_1 _12461_ (.CLK(clknet_leaf_81_mclk),
    .GATE(_00250_),
    .GCLK(_04486_));
 sky130_fd_sc_hd__dlclkp_1 _12462_ (.CLK(clknet_leaf_120_mclk),
    .GATE(net719),
    .GCLK(_04487_));
 sky130_fd_sc_hd__dlclkp_1 _12463_ (.CLK(clknet_leaf_117_mclk),
    .GATE(net719),
    .GCLK(_04488_));
 sky130_fd_sc_hd__dlclkp_1 _12464_ (.CLK(clknet_leaf_107_mclk),
    .GATE(net719),
    .GCLK(_04489_));
 sky130_fd_sc_hd__dlclkp_1 _12465_ (.CLK(clknet_leaf_90_mclk),
    .GATE(net721),
    .GCLK(_04490_));
 sky130_fd_sc_hd__dlclkp_1 _12466_ (.CLK(clknet_leaf_15_mclk),
    .GATE(net722),
    .GCLK(_04491_));
 sky130_fd_sc_hd__dlclkp_1 _12467_ (.CLK(clknet_leaf_107_mclk),
    .GATE(net721),
    .GCLK(_04492_));
 sky130_fd_sc_hd__dlclkp_4 _12468_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00251_),
    .GCLK(_04493_));
 sky130_fd_sc_hd__dlclkp_2 _12469_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00252_),
    .GCLK(_04494_));
 sky130_fd_sc_hd__dlclkp_2 _12470_ (.CLK(clknet_leaf_107_mclk),
    .GATE(_00253_),
    .GCLK(_04495_));
 sky130_fd_sc_hd__dlclkp_2 _12471_ (.CLK(clknet_leaf_105_mclk),
    .GATE(_00254_),
    .GCLK(_04496_));
 sky130_fd_sc_hd__dlclkp_2 _12472_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00255_),
    .GCLK(_04497_));
 sky130_fd_sc_hd__dlclkp_2 _12473_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00256_),
    .GCLK(_04498_));
 sky130_fd_sc_hd__dlclkp_2 _12474_ (.CLK(clknet_leaf_109_mclk),
    .GATE(_00257_),
    .GCLK(_04499_));
 sky130_fd_sc_hd__dlclkp_2 _12475_ (.CLK(clknet_leaf_106_mclk),
    .GATE(_00258_),
    .GCLK(_04500_));
 sky130_fd_sc_hd__dlclkp_2 _12476_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00259_),
    .GCLK(_04501_));
 sky130_fd_sc_hd__dlclkp_2 _12477_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00260_),
    .GCLK(_04502_));
 sky130_fd_sc_hd__dlclkp_2 _12478_ (.CLK(clknet_leaf_110_mclk),
    .GATE(_00261_),
    .GCLK(_04503_));
 sky130_fd_sc_hd__dlclkp_2 _12479_ (.CLK(clknet_leaf_104_mclk),
    .GATE(_00262_),
    .GCLK(_04504_));
 sky130_fd_sc_hd__dlclkp_2 _12480_ (.CLK(clknet_leaf_12_mclk),
    .GATE(_00263_),
    .GCLK(_04505_));
 sky130_fd_sc_hd__dlclkp_1 _12481_ (.CLK(clknet_leaf_80_mclk),
    .GATE(_00264_),
    .GCLK(_04506_));
 sky130_fd_sc_hd__dlclkp_1 _12482_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00265_),
    .GCLK(_04507_));
 sky130_fd_sc_hd__dlclkp_1 _12483_ (.CLK(clknet_leaf_12_mclk),
    .GATE(_00266_),
    .GCLK(_04508_));
 sky130_fd_sc_hd__dlclkp_1 _12484_ (.CLK(clknet_leaf_15_mclk),
    .GATE(_00267_),
    .GCLK(_04509_));
 sky130_fd_sc_hd__dlclkp_1 _12485_ (.CLK(clknet_leaf_13_mclk),
    .GATE(_00268_),
    .GCLK(_04510_));
 sky130_fd_sc_hd__dlclkp_1 _12486_ (.CLK(clknet_leaf_14_mclk),
    .GATE(_00269_),
    .GCLK(_04511_));
 sky130_fd_sc_hd__dlclkp_1 _12487_ (.CLK(clknet_leaf_19_mclk),
    .GATE(_00270_),
    .GCLK(_04512_));
 sky130_fd_sc_hd__dlclkp_1 _12488_ (.CLK(clknet_4_9__leaf_mclk),
    .GATE(_00271_),
    .GCLK(_04513_));
 sky130_fd_sc_hd__dlclkp_1 _12489_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00272_),
    .GCLK(_04514_));
 sky130_fd_sc_hd__dlclkp_1 _12490_ (.CLK(clknet_leaf_19_mclk),
    .GATE(_00273_),
    .GCLK(_04515_));
 sky130_fd_sc_hd__dlclkp_1 _12491_ (.CLK(clknet_leaf_22_mclk),
    .GATE(_00274_),
    .GCLK(_04516_));
 sky130_fd_sc_hd__dlclkp_1 _12492_ (.CLK(clknet_leaf_104_mclk),
    .GATE(_00275_),
    .GCLK(_04517_));
 sky130_fd_sc_hd__dlclkp_1 _12493_ (.CLK(clknet_leaf_20_mclk),
    .GATE(_00276_),
    .GCLK(_04518_));
 sky130_fd_sc_hd__dlclkp_1 _12494_ (.CLK(clknet_leaf_22_mclk),
    .GATE(_00277_),
    .GCLK(_04519_));
 sky130_fd_sc_hd__dlclkp_1 _12495_ (.CLK(clknet_leaf_17_mclk),
    .GATE(_00278_),
    .GCLK(_04520_));
 sky130_fd_sc_hd__dlclkp_1 _12496_ (.CLK(clknet_leaf_19_mclk),
    .GATE(_00279_),
    .GCLK(_04521_));
 sky130_fd_sc_hd__dlclkp_1 _12497_ (.CLK(clknet_leaf_112_mclk),
    .GATE(_00280_),
    .GCLK(_04522_));
 sky130_fd_sc_hd__dlclkp_1 _12498_ (.CLK(clknet_leaf_113_mclk),
    .GATE(_00281_),
    .GCLK(_04523_));
 sky130_fd_sc_hd__dlclkp_1 _12499_ (.CLK(clknet_leaf_114_mclk),
    .GATE(_00282_),
    .GCLK(_04524_));
 sky130_fd_sc_hd__dlclkp_1 _12500_ (.CLK(clknet_leaf_113_mclk),
    .GATE(_00283_),
    .GCLK(_04525_));
 sky130_fd_sc_hd__dlclkp_1 _12501_ (.CLK(clknet_leaf_109_mclk),
    .GATE(_00284_),
    .GCLK(_04526_));
 sky130_fd_sc_hd__dlclkp_1 _12502_ (.CLK(clknet_leaf_112_mclk),
    .GATE(_00285_),
    .GCLK(_04527_));
 sky130_fd_sc_hd__dlclkp_1 _12503_ (.CLK(clknet_leaf_80_mclk),
    .GATE(_00286_),
    .GCLK(_04528_));
 sky130_fd_sc_hd__dlclkp_1 _12504_ (.CLK(clknet_leaf_112_mclk),
    .GATE(_00287_),
    .GCLK(_04529_));
 sky130_fd_sc_hd__dlclkp_1 _12505_ (.CLK(clknet_leaf_113_mclk),
    .GATE(_00288_),
    .GCLK(_04530_));
 sky130_fd_sc_hd__dlclkp_1 _12506_ (.CLK(clknet_leaf_106_mclk),
    .GATE(_00289_),
    .GCLK(_04531_));
 sky130_fd_sc_hd__dlclkp_1 _12507_ (.CLK(clknet_leaf_105_mclk),
    .GATE(_00290_),
    .GCLK(_04532_));
 sky130_fd_sc_hd__dlclkp_1 _12508_ (.CLK(clknet_leaf_80_mclk),
    .GATE(_00291_),
    .GCLK(_04533_));
 sky130_fd_sc_hd__dlclkp_1 _12509_ (.CLK(clknet_leaf_106_mclk),
    .GATE(_00292_),
    .GCLK(_04534_));
 sky130_fd_sc_hd__dlclkp_1 _12510_ (.CLK(clknet_leaf_104_mclk),
    .GATE(_00293_),
    .GCLK(_04535_));
 sky130_fd_sc_hd__dlclkp_1 _12511_ (.CLK(clknet_leaf_16_mclk),
    .GATE(_00294_),
    .GCLK(_04536_));
 sky130_fd_sc_hd__dlclkp_1 _12512_ (.CLK(clknet_leaf_107_mclk),
    .GATE(_00295_),
    .GCLK(_04537_));
 sky130_fd_sc_hd__dlclkp_2 _12513_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00296_),
    .GCLK(_04538_));
 sky130_fd_sc_hd__dlclkp_2 _12514_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00297_),
    .GCLK(_04539_));
 sky130_fd_sc_hd__dlclkp_2 _12515_ (.CLK(clknet_leaf_80_mclk),
    .GATE(_00298_),
    .GCLK(_04540_));
 sky130_fd_sc_hd__dlclkp_2 _12516_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00299_),
    .GCLK(_04541_));
 sky130_fd_sc_hd__dlclkp_2 _12517_ (.CLK(clknet_leaf_21_mclk),
    .GATE(_00300_),
    .GCLK(_04542_));
 sky130_fd_sc_hd__dlclkp_2 _12518_ (.CLK(clknet_leaf_112_mclk),
    .GATE(_00301_),
    .GCLK(_04543_));
 sky130_fd_sc_hd__dlclkp_2 _12519_ (.CLK(clknet_leaf_106_mclk),
    .GATE(_00302_),
    .GCLK(_04544_));
 sky130_fd_sc_hd__dlclkp_2 _12520_ (.CLK(clknet_leaf_11_mclk),
    .GATE(_00303_),
    .GCLK(_04545_));
 sky130_fd_sc_hd__dlclkp_2 _12521_ (.CLK(clknet_leaf_53_mclk),
    .GATE(_00304_),
    .GCLK(_04546_));
 sky130_fd_sc_hd__dlclkp_2 _12522_ (.CLK(clknet_leaf_111_mclk),
    .GATE(_00305_),
    .GCLK(_04547_));
 sky130_fd_sc_hd__dlclkp_2 _12523_ (.CLK(clknet_4_6__leaf_mclk),
    .GATE(_00306_),
    .GCLK(_04548_));
 sky130_fd_sc_hd__dlclkp_2 _12524_ (.CLK(clknet_leaf_12_mclk),
    .GATE(_00307_),
    .GCLK(_04549_));
 sky130_fd_sc_hd__dlclkp_4 _12525_ (.CLK(clknet_leaf_79_mclk),
    .GATE(_00311_),
    .GCLK(_04550_));
 sky130_fd_sc_hd__dlclkp_1 _12526_ (.CLK(clknet_leaf_82_mclk),
    .GATE(_00312_),
    .GCLK(_04551_));
 sky130_fd_sc_hd__dlclkp_1 _12527_ (.CLK(clknet_leaf_81_mclk),
    .GATE(_00313_),
    .GCLK(_04552_));
 sky130_fd_sc_hd__dlclkp_1 _12528_ (.CLK(clknet_leaf_87_mclk),
    .GATE(_00314_),
    .GCLK(_04553_));
 sky130_fd_sc_hd__dlclkp_1 _12529_ (.CLK(clknet_leaf_87_mclk),
    .GATE(_00315_),
    .GCLK(_04554_));
 sky130_fd_sc_hd__dlclkp_1 _12530_ (.CLK(clknet_leaf_83_mclk),
    .GATE(_00316_),
    .GCLK(_04555_));
 sky130_fd_sc_hd__dlclkp_1 _12531_ (.CLK(clknet_leaf_87_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04556_));
 sky130_fd_sc_hd__dlclkp_1 _12532_ (.CLK(clknet_leaf_87_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04557_));
 sky130_fd_sc_hd__dlclkp_1 _12533_ (.CLK(clknet_leaf_83_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04558_));
 sky130_fd_sc_hd__dlclkp_1 _12534_ (.CLK(clknet_leaf_76_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04559_));
 sky130_fd_sc_hd__dlclkp_1 _12535_ (.CLK(clknet_leaf_76_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04560_));
 sky130_fd_sc_hd__dlclkp_1 _12536_ (.CLK(clknet_leaf_75_mclk),
    .GATE(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04561_));
 sky130_fd_sc_hd__dlclkp_2 _12537_ (.CLK(clknet_leaf_72_mclk),
    .GATE(_00350_),
    .GCLK(_04562_));
 sky130_fd_sc_hd__dlclkp_1 _12538_ (.CLK(clknet_leaf_78_mclk),
    .GATE(_00351_),
    .GCLK(_04563_));
 sky130_fd_sc_hd__dlclkp_4 _12539_ (.CLK(clknet_leaf_79_mclk),
    .GATE(_00352_),
    .GCLK(_04564_));
 sky130_fd_sc_hd__dlclkp_4 _12540_ (.CLK(clknet_leaf_76_mclk),
    .GATE(_00353_),
    .GCLK(_04565_));
 sky130_fd_sc_hd__dlclkp_4 _12541_ (.CLK(clknet_leaf_76_mclk),
    .GATE(_00353_),
    .GCLK(_04566_));
 sky130_fd_sc_hd__dlclkp_4 _12542_ (.CLK(clknet_leaf_76_mclk),
    .GATE(_00353_),
    .GCLK(_04567_));
 sky130_fd_sc_hd__dlclkp_2 _12543_ (.CLK(clknet_leaf_79_mclk),
    .GATE(_00354_),
    .GCLK(_04568_));
 sky130_fd_sc_hd__dlclkp_2 _12544_ (.CLK(clknet_leaf_58_mclk),
    .GATE(_00355_),
    .GCLK(_04569_));
 sky130_fd_sc_hd__dlclkp_2 _12545_ (.CLK(clknet_leaf_77_mclk),
    .GATE(_00356_),
    .GCLK(_04570_));
 sky130_fd_sc_hd__dlclkp_2 _12546_ (.CLK(clknet_leaf_78_mclk),
    .GATE(_00357_),
    .GCLK(_04571_));
 sky130_fd_sc_hd__dlclkp_2 _12547_ (.CLK(clknet_4_12__leaf_mclk),
    .GATE(_00358_),
    .GCLK(_04572_));
 sky130_fd_sc_hd__dlclkp_2 _12548_ (.CLK(clknet_leaf_60_mclk),
    .GATE(_00359_),
    .GCLK(_04573_));
 sky130_fd_sc_hd__dlclkp_2 _12549_ (.CLK(clknet_leaf_77_mclk),
    .GATE(_00360_),
    .GCLK(_04574_));
 sky130_fd_sc_hd__dlclkp_2 _12550_ (.CLK(clknet_leaf_78_mclk),
    .GATE(_00361_),
    .GCLK(_04575_));
 sky130_fd_sc_hd__dlclkp_2 _12551_ (.CLK(clknet_leaf_60_mclk),
    .GATE(_00362_),
    .GCLK(_04576_));
 sky130_fd_sc_hd__dlclkp_2 _12552_ (.CLK(clknet_leaf_60_mclk),
    .GATE(_00363_),
    .GCLK(_04577_));
 sky130_fd_sc_hd__dlclkp_2 _12553_ (.CLK(clknet_leaf_77_mclk),
    .GATE(_00364_),
    .GCLK(_04578_));
 sky130_fd_sc_hd__dlclkp_2 _12554_ (.CLK(clknet_leaf_78_mclk),
    .GATE(_00365_),
    .GCLK(_04579_));
 sky130_fd_sc_hd__dlclkp_2 _12555_ (.CLK(clknet_4_12__leaf_mclk),
    .GATE(_00366_),
    .GCLK(_04580_));
 sky130_fd_sc_hd__dlclkp_2 _12556_ (.CLK(clknet_leaf_60_mclk),
    .GATE(_00367_),
    .GCLK(_04581_));
 sky130_fd_sc_hd__dlclkp_2 _12557_ (.CLK(clknet_4_13__leaf_mclk),
    .GATE(_00368_),
    .GCLK(_04582_));
 sky130_fd_sc_hd__dlclkp_2 _12558_ (.CLK(clknet_leaf_78_mclk),
    .GATE(_00369_),
    .GCLK(_04583_));
 sky130_fd_sc_hd__dlclkp_2 _12559_ (.CLK(clknet_leaf_91_mclk),
    .GATE(_00403_),
    .GCLK(_04584_));
 sky130_fd_sc_hd__dlclkp_1 _12560_ (.CLK(clknet_leaf_84_mclk),
    .GATE(_00404_),
    .GCLK(_04585_));
 sky130_fd_sc_hd__dlclkp_4 _12561_ (.CLK(clknet_leaf_80_mclk),
    .GATE(_00405_),
    .GCLK(_04586_));
 sky130_fd_sc_hd__dlclkp_4 _12562_ (.CLK(clknet_leaf_87_mclk),
    .GATE(_00406_),
    .GCLK(_04587_));
 sky130_fd_sc_hd__dlclkp_4 _12563_ (.CLK(clknet_leaf_83_mclk),
    .GATE(_00406_),
    .GCLK(_04588_));
 sky130_fd_sc_hd__dlclkp_4 _12564_ (.CLK(clknet_leaf_86_mclk),
    .GATE(_00406_),
    .GCLK(_04589_));
 sky130_fd_sc_hd__dlclkp_2 _12565_ (.CLK(clknet_leaf_85_mclk),
    .GATE(_00407_),
    .GCLK(_04590_));
 sky130_fd_sc_hd__dlclkp_2 _12566_ (.CLK(clknet_leaf_102_mclk),
    .GATE(_00408_),
    .GCLK(_04591_));
 sky130_fd_sc_hd__dlclkp_2 _12567_ (.CLK(clknet_leaf_86_mclk),
    .GATE(_00409_),
    .GCLK(_04592_));
 sky130_fd_sc_hd__dlclkp_2 _12568_ (.CLK(clknet_leaf_82_mclk),
    .GATE(_00410_),
    .GCLK(_04593_));
 sky130_fd_sc_hd__dlclkp_2 _12569_ (.CLK(clknet_leaf_85_mclk),
    .GATE(_00411_),
    .GCLK(_04594_));
 sky130_fd_sc_hd__dlclkp_2 _12570_ (.CLK(clknet_leaf_105_mclk),
    .GATE(_00412_),
    .GCLK(_04595_));
 sky130_fd_sc_hd__dlclkp_2 _12571_ (.CLK(clknet_leaf_86_mclk),
    .GATE(_00413_),
    .GCLK(_04596_));
 sky130_fd_sc_hd__dlclkp_2 _12572_ (.CLK(clknet_leaf_84_mclk),
    .GATE(_00414_),
    .GCLK(_04597_));
 sky130_fd_sc_hd__dlclkp_2 _12573_ (.CLK(clknet_4_4__leaf_mclk),
    .GATE(_00415_),
    .GCLK(_04598_));
 sky130_fd_sc_hd__dlclkp_2 _12574_ (.CLK(clknet_leaf_103_mclk),
    .GATE(_00416_),
    .GCLK(_04599_));
 sky130_fd_sc_hd__dlclkp_2 _12575_ (.CLK(clknet_leaf_86_mclk),
    .GATE(_00417_),
    .GCLK(_04600_));
 sky130_fd_sc_hd__dlclkp_2 _12576_ (.CLK(clknet_leaf_84_mclk),
    .GATE(_00418_),
    .GCLK(_04601_));
 sky130_fd_sc_hd__dlclkp_2 _12577_ (.CLK(clknet_leaf_85_mclk),
    .GATE(_00419_),
    .GCLK(_04602_));
 sky130_fd_sc_hd__dlclkp_2 _12578_ (.CLK(clknet_leaf_102_mclk),
    .GATE(_00420_),
    .GCLK(_04603_));
 sky130_fd_sc_hd__dlclkp_2 _12579_ (.CLK(clknet_leaf_86_mclk),
    .GATE(_00421_),
    .GCLK(_04604_));
 sky130_fd_sc_hd__dlclkp_2 _12580_ (.CLK(clknet_leaf_84_mclk),
    .GATE(_00422_),
    .GCLK(_04605_));
 sky130_fd_sc_hd__dlclkp_2 _12581_ (.CLK(clknet_leaf_94_mclk),
    .GATE(_00456_),
    .GCLK(_04606_));
 sky130_fd_sc_hd__dlclkp_1 _12582_ (.CLK(clknet_leaf_103_mclk),
    .GATE(_00457_),
    .GCLK(_04607_));
 sky130_fd_sc_hd__dlclkp_4 _12583_ (.CLK(clknet_leaf_103_mclk),
    .GATE(_00458_),
    .GCLK(_04608_));
 sky130_fd_sc_hd__dlclkp_4 _12584_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00459_),
    .GCLK(_04609_));
 sky130_fd_sc_hd__dlclkp_4 _12585_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00459_),
    .GCLK(_04610_));
 sky130_fd_sc_hd__dlclkp_4 _12586_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00459_),
    .GCLK(_04611_));
 sky130_fd_sc_hd__dlclkp_2 _12587_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00460_),
    .GCLK(_04612_));
 sky130_fd_sc_hd__dlclkp_2 _12588_ (.CLK(clknet_leaf_114_mclk),
    .GATE(_00461_),
    .GCLK(_04613_));
 sky130_fd_sc_hd__dlclkp_2 _12589_ (.CLK(clknet_leaf_96_mclk),
    .GATE(_00462_),
    .GCLK(_04614_));
 sky130_fd_sc_hd__dlclkp_2 _12590_ (.CLK(clknet_leaf_99_mclk),
    .GATE(_00463_),
    .GCLK(_04615_));
 sky130_fd_sc_hd__dlclkp_2 _12591_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00464_),
    .GCLK(_04616_));
 sky130_fd_sc_hd__dlclkp_2 _12592_ (.CLK(clknet_leaf_115_mclk),
    .GATE(_00465_),
    .GCLK(_04617_));
 sky130_fd_sc_hd__dlclkp_2 _12593_ (.CLK(clknet_leaf_97_mclk),
    .GATE(_00466_),
    .GCLK(_04618_));
 sky130_fd_sc_hd__dlclkp_2 _12594_ (.CLK(clknet_leaf_99_mclk),
    .GATE(_00467_),
    .GCLK(_04619_));
 sky130_fd_sc_hd__dlclkp_2 _12595_ (.CLK(clknet_leaf_100_mclk),
    .GATE(_00468_),
    .GCLK(_04620_));
 sky130_fd_sc_hd__dlclkp_2 _12596_ (.CLK(clknet_leaf_116_mclk),
    .GATE(_00469_),
    .GCLK(_04621_));
 sky130_fd_sc_hd__dlclkp_2 _12597_ (.CLK(clknet_leaf_96_mclk),
    .GATE(_00470_),
    .GCLK(_04622_));
 sky130_fd_sc_hd__dlclkp_2 _12598_ (.CLK(clknet_leaf_99_mclk),
    .GATE(_00471_),
    .GCLK(_04623_));
 sky130_fd_sc_hd__dlclkp_2 _12599_ (.CLK(clknet_leaf_97_mclk),
    .GATE(_00472_),
    .GCLK(_04624_));
 sky130_fd_sc_hd__dlclkp_2 _12600_ (.CLK(clknet_leaf_116_mclk),
    .GATE(_00473_),
    .GCLK(_04625_));
 sky130_fd_sc_hd__dlclkp_2 _12601_ (.CLK(clknet_4_5__leaf_mclk),
    .GATE(_00474_),
    .GCLK(_04626_));
 sky130_fd_sc_hd__dlclkp_2 _12602_ (.CLK(clknet_leaf_99_mclk),
    .GATE(_00475_),
    .GCLK(_04627_));
 sky130_fd_sc_hd__dlclkp_2 _12603_ (.CLK(clknet_leaf_55_mclk),
    .GATE(_00476_),
    .GCLK(_04628_));
 sky130_fd_sc_hd__dlclkp_2 _12604_ (.CLK(clknet_leaf_55_mclk),
    .GATE(_00477_),
    .GCLK(_04629_));
 sky130_fd_sc_hd__dlclkp_2 _12605_ (.CLK(clknet_leaf_58_mclk),
    .GATE(_00478_),
    .GCLK(_04630_));
 sky130_fd_sc_hd__dlclkp_2 _12606_ (.CLK(clknet_leaf_46_mclk),
    .GATE(\u_gpio.pulse_1us ),
    .GCLK(_04631_));
 sky130_fd_sc_hd__dlclkp_2 _12607_ (.CLK(clknet_leaf_117_mclk),
    .GATE(net533),
    .GCLK(_04632_));
 sky130_fd_sc_hd__dlclkp_4 _12608_ (.CLK(clknet_leaf_55_mclk),
    .GATE(_00510_),
    .GCLK(_04633_));
 sky130_fd_sc_hd__dlclkp_2 _12609_ (.CLK(clknet_leaf_54_mclk),
    .GATE(_00511_),
    .GCLK(_04634_));
 sky130_fd_sc_hd__dlclkp_2 _12610_ (.CLK(clknet_leaf_17_mclk),
    .GATE(_00512_),
    .GCLK(_04635_));
 sky130_fd_sc_hd__dlclkp_2 _12611_ (.CLK(clknet_leaf_47_mclk),
    .GATE(_00513_),
    .GCLK(_04636_));
 sky130_fd_sc_hd__dlclkp_2 _12612_ (.CLK(clknet_leaf_51_mclk),
    .GATE(_00514_),
    .GCLK(_04637_));
 sky130_fd_sc_hd__dlclkp_2 _12613_ (.CLK(clknet_leaf_51_mclk),
    .GATE(_00515_),
    .GCLK(_04638_));
 sky130_fd_sc_hd__dlclkp_2 _12614_ (.CLK(clknet_leaf_17_mclk),
    .GATE(_00516_),
    .GCLK(_04639_));
 sky130_fd_sc_hd__dlclkp_2 _12615_ (.CLK(clknet_4_11__leaf_mclk),
    .GATE(_00517_),
    .GCLK(_04640_));
 sky130_fd_sc_hd__dlclkp_2 _12616_ (.CLK(clknet_leaf_51_mclk),
    .GATE(_00518_),
    .GCLK(_04641_));
 sky130_fd_sc_hd__dlclkp_2 _12617_ (.CLK(clknet_leaf_53_mclk),
    .GATE(_00519_),
    .GCLK(_04642_));
 sky130_fd_sc_hd__dlclkp_2 _12618_ (.CLK(clknet_leaf_17_mclk),
    .GATE(_00520_),
    .GCLK(_04643_));
 sky130_fd_sc_hd__dlclkp_2 _12619_ (.CLK(clknet_leaf_45_mclk),
    .GATE(_00521_),
    .GCLK(_04644_));
 sky130_fd_sc_hd__dlclkp_2 _12620_ (.CLK(clknet_4_11__leaf_mclk),
    .GATE(_00522_),
    .GCLK(_04645_));
 sky130_fd_sc_hd__dlclkp_2 _12621_ (.CLK(clknet_leaf_53_mclk),
    .GATE(_00523_),
    .GCLK(_04646_));
 sky130_fd_sc_hd__dlclkp_2 _12622_ (.CLK(clknet_leaf_17_mclk),
    .GATE(_00524_),
    .GCLK(_04647_));
 sky130_fd_sc_hd__dlclkp_2 _12623_ (.CLK(clknet_leaf_45_mclk),
    .GATE(_00525_),
    .GCLK(_04648_));
 sky130_fd_sc_hd__dlclkp_2 _12624_ (.CLK(clknet_leaf_45_mclk),
    .GATE(_00526_),
    .GCLK(_04649_));
 sky130_fd_sc_hd__dlclkp_2 _12625_ (.CLK(clknet_leaf_54_mclk),
    .GATE(_00543_),
    .GCLK(_04650_));
 sky130_fd_sc_hd__dlclkp_2 _12626_ (.CLK(clknet_leaf_53_mclk),
    .GATE(_00560_),
    .GCLK(_04651_));
 sky130_fd_sc_hd__dlclkp_2 _12627_ (.CLK(clknet_leaf_53_mclk),
    .GATE(_00577_),
    .GCLK(_04652_));
 sky130_fd_sc_hd__dlclkp_4 _12628_ (.CLK(clknet_leaf_63_mclk),
    .GATE(_00579_),
    .GCLK(_04653_));
 sky130_fd_sc_hd__dlclkp_1 _12629_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00582_),
    .GCLK(_04654_));
 sky130_fd_sc_hd__dlclkp_1 _12630_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00583_),
    .GCLK(_04655_));
 sky130_fd_sc_hd__dlclkp_1 _12631_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00584_),
    .GCLK(_04656_));
 sky130_fd_sc_hd__dlclkp_1 _12632_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00584_),
    .GCLK(_04657_));
 sky130_fd_sc_hd__dlclkp_4 _12633_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00585_),
    .GCLK(_04658_));
 sky130_fd_sc_hd__dlclkp_4 _12634_ (.CLK(clknet_leaf_62_mclk),
    .GATE(_00586_),
    .GCLK(_04659_));
 sky130_fd_sc_hd__dlclkp_1 _12635_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00589_),
    .GCLK(_04660_));
 sky130_fd_sc_hd__dlclkp_1 _12636_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00590_),
    .GCLK(_04661_));
 sky130_fd_sc_hd__dlclkp_1 _12637_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00591_),
    .GCLK(_04662_));
 sky130_fd_sc_hd__dlclkp_1 _12638_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00591_),
    .GCLK(_04663_));
 sky130_fd_sc_hd__dlclkp_4 _12639_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00592_),
    .GCLK(_04664_));
 sky130_fd_sc_hd__dlclkp_4 _12640_ (.CLK(clknet_leaf_66_mclk),
    .GATE(_00593_),
    .GCLK(_04665_));
 sky130_fd_sc_hd__dlclkp_1 _12641_ (.CLK(clknet_leaf_67_mclk),
    .GATE(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04666_));
 sky130_fd_sc_hd__dlclkp_1 _12642_ (.CLK(clknet_leaf_67_mclk),
    .GATE(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04667_));
 sky130_fd_sc_hd__dlclkp_1 _12643_ (.CLK(clknet_leaf_67_mclk),
    .GATE(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04668_));
 sky130_fd_sc_hd__dlclkp_1 _12644_ (.CLK(clknet_leaf_62_mclk),
    .GATE(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[0].u_bit_reg.we ),
    .GCLK(_04669_));
 sky130_fd_sc_hd__dlclkp_2 _12645_ (.CLK(clknet_4_14__leaf_mclk),
    .GATE(_00594_),
    .GCLK(_04670_));
 sky130_fd_sc_hd__dlclkp_2 _12646_ (.CLK(clknet_leaf_67_mclk),
    .GATE(_00595_),
    .GCLK(_04671_));
 sky130_fd_sc_hd__dlclkp_2 _12647_ (.CLK(clknet_leaf_65_mclk),
    .GATE(_00596_),
    .GCLK(_04672_));
 sky130_fd_sc_hd__dlclkp_2 _12648_ (.CLK(clknet_4_14__leaf_mclk),
    .GATE(_00597_),
    .GCLK(_04673_));
 sky130_fd_sc_hd__dlclkp_2 _12649_ (.CLK(clknet_leaf_67_mclk),
    .GATE(_00598_),
    .GCLK(_04674_));
 sky130_fd_sc_hd__dlclkp_2 _12650_ (.CLK(clknet_leaf_65_mclk),
    .GATE(_00599_),
    .GCLK(_04675_));
 sky130_fd_sc_hd__dlclkp_2 _12651_ (.CLK(clknet_leaf_70_mclk),
    .GATE(_00647_),
    .GCLK(_04676_));
 sky130_fd_sc_hd__dlclkp_1 _12652_ (.CLK(clknet_leaf_70_mclk),
    .GATE(_00648_),
    .GCLK(_04677_));
 sky130_fd_sc_hd__dlclkp_1 _12653_ (.CLK(clknet_leaf_67_mclk),
    .GATE(_00649_),
    .GCLK(_04678_));
 sky130_fd_sc_hd__dlclkp_2 _12654_ (.CLK(clknet_4_15__leaf_mclk),
    .GATE(_00650_),
    .GCLK(_04679_));
 sky130_fd_sc_hd__dlclkp_4 _12655_ (.CLK(clknet_leaf_67_mclk),
    .GATE(_00647_),
    .GCLK(_04680_));
 sky130_fd_sc_hd__dlclkp_2 _12656_ (.CLK(clknet_leaf_69_mclk),
    .GATE(_00698_),
    .GCLK(_04682_));
 sky130_fd_sc_hd__dlclkp_1 _12657_ (.CLK(clknet_leaf_69_mclk),
    .GATE(_00699_),
    .GCLK(_04683_));
 sky130_fd_sc_hd__dlclkp_1 _12658_ (.CLK(clknet_leaf_69_mclk),
    .GATE(_00700_),
    .GCLK(_04684_));
 sky130_fd_sc_hd__dlclkp_2 _12659_ (.CLK(clknet_leaf_69_mclk),
    .GATE(_00701_),
    .GCLK(_04685_));
 sky130_fd_sc_hd__dlclkp_4 _12660_ (.CLK(clknet_leaf_69_mclk),
    .GATE(_00698_),
    .GCLK(_04686_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04347_ (.A(_04347_),
    .X(clknet_0__04347_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04353_ (.A(_04353_),
    .X(clknet_0__04353_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04354_ (.A(_04354_),
    .X(clknet_0__04354_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04355_ (.A(_04355_),
    .X(clknet_0__04355_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04356_ (.A(_04356_),
    .X(clknet_0__04356_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04357_ (.A(_04357_),
    .X(clknet_0__04357_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04358_ (.A(_04358_),
    .X(clknet_0__04358_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04359_ (.A(_04359_),
    .X(clknet_0__04359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04392_ (.A(_04392_),
    .X(clknet_0__04392_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04393_ (.A(_04393_),
    .X(clknet_0__04393_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04394_ (.A(_04394_),
    .X(clknet_0__04394_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04395_ (.A(_04395_),
    .X(clknet_0__04395_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04396_ (.A(_04396_),
    .X(clknet_0__04396_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04397_ (.A(_04397_),
    .X(clknet_0__04397_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04398_ (.A(_04398_),
    .X(clknet_0__04398_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04399_ (.A(_04399_),
    .X(clknet_0__04399_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04400_ (.A(_04400_),
    .X(clknet_0__04400_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04401_ (.A(_04401_),
    .X(clknet_0__04401_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04402_ (.A(_04402_),
    .X(clknet_0__04402_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04403_ (.A(_04403_),
    .X(clknet_0__04403_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04404_ (.A(_04404_),
    .X(clknet_0__04404_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04405_ (.A(_04405_),
    .X(clknet_0__04405_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04406_ (.A(_04406_),
    .X(clknet_0__04406_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04407_ (.A(_04407_),
    .X(clknet_0__04407_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04408_ (.A(_04408_),
    .X(clknet_0__04408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04409_ (.A(_04409_),
    .X(clknet_0__04409_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04410_ (.A(_04410_),
    .X(clknet_0__04410_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04411_ (.A(_04411_),
    .X(clknet_0__04411_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04412_ (.A(_04412_),
    .X(clknet_0__04412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04413_ (.A(_04413_),
    .X(clknet_0__04413_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04414_ (.A(_04414_),
    .X(clknet_0__04414_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04415_ (.A(_04415_),
    .X(clknet_0__04415_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04416_ (.A(_04416_),
    .X(clknet_0__04416_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04417_ (.A(_04417_),
    .X(clknet_0__04417_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04418_ (.A(_04418_),
    .X(clknet_0__04418_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04419_ (.A(_04419_),
    .X(clknet_0__04419_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04420_ (.A(_04420_),
    .X(clknet_0__04420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04421_ (.A(_04421_),
    .X(clknet_0__04421_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04422_ (.A(_04422_),
    .X(clknet_0__04422_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04423_ (.A(_04423_),
    .X(clknet_0__04423_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04424_ (.A(_04424_),
    .X(clknet_0__04424_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04425_ (.A(_04425_),
    .X(clknet_0__04425_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04426_ (.A(_04426_),
    .X(clknet_0__04426_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04427_ (.A(_04427_),
    .X(clknet_0__04427_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04428_ (.A(_04428_),
    .X(clknet_0__04428_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04429_ (.A(_04429_),
    .X(clknet_0__04429_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04430_ (.A(_04430_),
    .X(clknet_0__04430_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04431_ (.A(_04431_),
    .X(clknet_0__04431_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04432_ (.A(_04432_),
    .X(clknet_0__04432_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04433_ (.A(_04433_),
    .X(clknet_0__04433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04434_ (.A(_04434_),
    .X(clknet_0__04434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04435_ (.A(_04435_),
    .X(clknet_0__04435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04436_ (.A(_04436_),
    .X(clknet_0__04436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04437_ (.A(_04437_),
    .X(clknet_0__04437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04438_ (.A(_04438_),
    .X(clknet_0__04438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04439_ (.A(_04439_),
    .X(clknet_0__04439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04440_ (.A(_04440_),
    .X(clknet_0__04440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04441_ (.A(_04441_),
    .X(clknet_0__04441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04442_ (.A(_04442_),
    .X(clknet_0__04442_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04443_ (.A(_04443_),
    .X(clknet_0__04443_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04444_ (.A(_04444_),
    .X(clknet_0__04444_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04445_ (.A(_04445_),
    .X(clknet_0__04445_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04446_ (.A(_04446_),
    .X(clknet_0__04446_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04447_ (.A(_04447_),
    .X(clknet_0__04447_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04448_ (.A(_04448_),
    .X(clknet_0__04448_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04449_ (.A(_04449_),
    .X(clknet_0__04449_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04450_ (.A(_04450_),
    .X(clknet_0__04450_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04451_ (.A(_04451_),
    .X(clknet_0__04451_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04452_ (.A(_04452_),
    .X(clknet_0__04452_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04453_ (.A(_04453_),
    .X(clknet_0__04453_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04454_ (.A(_04454_),
    .X(clknet_0__04454_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04455_ (.A(_04455_),
    .X(clknet_0__04455_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04456_ (.A(_04456_),
    .X(clknet_0__04456_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04457_ (.A(_04457_),
    .X(clknet_0__04457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04458_ (.A(_04458_),
    .X(clknet_0__04458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04459_ (.A(_04459_),
    .X(clknet_0__04459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04460_ (.A(_04460_),
    .X(clknet_0__04460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04461_ (.A(_04461_),
    .X(clknet_0__04461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04463_ (.A(_04463_),
    .X(clknet_0__04463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04464_ (.A(_04464_),
    .X(clknet_0__04464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04465_ (.A(_04465_),
    .X(clknet_0__04465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04466_ (.A(_04466_),
    .X(clknet_0__04466_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04467_ (.A(_04467_),
    .X(clknet_0__04467_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04468_ (.A(_04468_),
    .X(clknet_0__04468_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04469_ (.A(_04469_),
    .X(clknet_0__04469_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04470_ (.A(_04470_),
    .X(clknet_0__04470_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04471_ (.A(_04471_),
    .X(clknet_0__04471_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04472_ (.A(_04472_),
    .X(clknet_0__04472_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04473_ (.A(_04473_),
    .X(clknet_0__04473_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04474_ (.A(_04474_),
    .X(clknet_0__04474_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04475_ (.A(_04475_),
    .X(clknet_0__04475_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04476_ (.A(_04476_),
    .X(clknet_0__04476_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04477_ (.A(_04477_),
    .X(clknet_0__04477_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04478_ (.A(_04478_),
    .X(clknet_0__04478_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04479_ (.A(_04479_),
    .X(clknet_0__04479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04480_ (.A(_04480_),
    .X(clknet_0__04480_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04481_ (.A(_04481_),
    .X(clknet_0__04481_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04482_ (.A(_04482_),
    .X(clknet_0__04482_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04483_ (.A(_04483_),
    .X(clknet_0__04483_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04484_ (.A(_04484_),
    .X(clknet_0__04484_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04485_ (.A(_04485_),
    .X(clknet_0__04485_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04486_ (.A(_04486_),
    .X(clknet_0__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04487_ (.A(_04487_),
    .X(clknet_0__04487_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04488_ (.A(_04488_),
    .X(clknet_0__04488_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04489_ (.A(_04489_),
    .X(clknet_0__04489_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04490_ (.A(_04490_),
    .X(clknet_0__04490_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04491_ (.A(_04491_),
    .X(clknet_0__04491_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04492_ (.A(_04492_),
    .X(clknet_0__04492_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04493_ (.A(_04493_),
    .X(clknet_0__04493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04494_ (.A(_04494_),
    .X(clknet_0__04494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04495_ (.A(_04495_),
    .X(clknet_0__04495_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04496_ (.A(_04496_),
    .X(clknet_0__04496_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04497_ (.A(_04497_),
    .X(clknet_0__04497_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04498_ (.A(_04498_),
    .X(clknet_0__04498_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04499_ (.A(_04499_),
    .X(clknet_0__04499_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04500_ (.A(_04500_),
    .X(clknet_0__04500_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04501_ (.A(_04501_),
    .X(clknet_0__04501_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04502_ (.A(_04502_),
    .X(clknet_0__04502_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04503_ (.A(_04503_),
    .X(clknet_0__04503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04504_ (.A(_04504_),
    .X(clknet_0__04504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04505_ (.A(_04505_),
    .X(clknet_0__04505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04538_ (.A(_04538_),
    .X(clknet_0__04538_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04539_ (.A(_04539_),
    .X(clknet_0__04539_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04540_ (.A(_04540_),
    .X(clknet_0__04540_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04541_ (.A(_04541_),
    .X(clknet_0__04541_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04542_ (.A(_04542_),
    .X(clknet_0__04542_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04543_ (.A(_04543_),
    .X(clknet_0__04543_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04544_ (.A(_04544_),
    .X(clknet_0__04544_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04545_ (.A(_04545_),
    .X(clknet_0__04545_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04546_ (.A(_04546_),
    .X(clknet_0__04546_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04547_ (.A(_04547_),
    .X(clknet_0__04547_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04548_ (.A(_04548_),
    .X(clknet_0__04548_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04549_ (.A(_04549_),
    .X(clknet_0__04549_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04550_ (.A(_04550_),
    .X(clknet_0__04550_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04551_ (.A(_04551_),
    .X(clknet_0__04551_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04552_ (.A(_04552_),
    .X(clknet_0__04552_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04562_ (.A(_04562_),
    .X(clknet_0__04562_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04564_ (.A(_04564_),
    .X(clknet_0__04564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04565_ (.A(_04565_),
    .X(clknet_0__04565_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04566_ (.A(_04566_),
    .X(clknet_0__04566_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04567_ (.A(_04567_),
    .X(clknet_0__04567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04568_ (.A(_04568_),
    .X(clknet_0__04568_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04569_ (.A(_04569_),
    .X(clknet_0__04569_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04570_ (.A(_04570_),
    .X(clknet_0__04570_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04571_ (.A(_04571_),
    .X(clknet_0__04571_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04572_ (.A(_04572_),
    .X(clknet_0__04572_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04573_ (.A(_04573_),
    .X(clknet_0__04573_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04574_ (.A(_04574_),
    .X(clknet_0__04574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04575_ (.A(_04575_),
    .X(clknet_0__04575_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04576_ (.A(_04576_),
    .X(clknet_0__04576_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04577_ (.A(_04577_),
    .X(clknet_0__04577_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04578_ (.A(_04578_),
    .X(clknet_0__04578_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04579_ (.A(_04579_),
    .X(clknet_0__04579_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04580_ (.A(_04580_),
    .X(clknet_0__04580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04581_ (.A(_04581_),
    .X(clknet_0__04581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04582_ (.A(_04582_),
    .X(clknet_0__04582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04583_ (.A(_04583_),
    .X(clknet_0__04583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04584_ (.A(_04584_),
    .X(clknet_0__04584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04586_ (.A(_04586_),
    .X(clknet_0__04586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04587_ (.A(_04587_),
    .X(clknet_0__04587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04588_ (.A(_04588_),
    .X(clknet_0__04588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04589_ (.A(_04589_),
    .X(clknet_0__04589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04590_ (.A(_04590_),
    .X(clknet_0__04590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04591_ (.A(_04591_),
    .X(clknet_0__04591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04592_ (.A(_04592_),
    .X(clknet_0__04592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04593_ (.A(_04593_),
    .X(clknet_0__04593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04594_ (.A(_04594_),
    .X(clknet_0__04594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04595_ (.A(_04595_),
    .X(clknet_0__04595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04596_ (.A(_04596_),
    .X(clknet_0__04596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04597_ (.A(_04597_),
    .X(clknet_0__04597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04598_ (.A(_04598_),
    .X(clknet_0__04598_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04599_ (.A(_04599_),
    .X(clknet_0__04599_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04600_ (.A(_04600_),
    .X(clknet_0__04600_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04601_ (.A(_04601_),
    .X(clknet_0__04601_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04602_ (.A(_04602_),
    .X(clknet_0__04602_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04603_ (.A(_04603_),
    .X(clknet_0__04603_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04604_ (.A(_04604_),
    .X(clknet_0__04604_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04605_ (.A(_04605_),
    .X(clknet_0__04605_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04606_ (.A(_04606_),
    .X(clknet_0__04606_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04608_ (.A(_04608_),
    .X(clknet_0__04608_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04609_ (.A(_04609_),
    .X(clknet_0__04609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04610_ (.A(_04610_),
    .X(clknet_0__04610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04611_ (.A(_04611_),
    .X(clknet_0__04611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04612_ (.A(_04612_),
    .X(clknet_0__04612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04613_ (.A(_04613_),
    .X(clknet_0__04613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04614_ (.A(_04614_),
    .X(clknet_0__04614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04615_ (.A(_04615_),
    .X(clknet_0__04615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04616_ (.A(_04616_),
    .X(clknet_0__04616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04617_ (.A(_04617_),
    .X(clknet_0__04617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04618_ (.A(_04618_),
    .X(clknet_0__04618_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04619_ (.A(_04619_),
    .X(clknet_0__04619_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04620_ (.A(_04620_),
    .X(clknet_0__04620_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04621_ (.A(_04621_),
    .X(clknet_0__04621_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04622_ (.A(_04622_),
    .X(clknet_0__04622_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04623_ (.A(_04623_),
    .X(clknet_0__04623_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04624_ (.A(_04624_),
    .X(clknet_0__04624_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04625_ (.A(_04625_),
    .X(clknet_0__04625_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04626_ (.A(_04626_),
    .X(clknet_0__04626_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04627_ (.A(_04627_),
    .X(clknet_0__04627_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04628_ (.A(_04628_),
    .X(clknet_0__04628_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04629_ (.A(_04629_),
    .X(clknet_0__04629_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04630_ (.A(_04630_),
    .X(clknet_0__04630_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04631_ (.A(_04631_),
    .X(clknet_0__04631_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04632_ (.A(_04632_),
    .X(clknet_0__04632_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04633_ (.A(_04633_),
    .X(clknet_0__04633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04634_ (.A(_04634_),
    .X(clknet_0__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04635_ (.A(_04635_),
    .X(clknet_0__04635_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04636_ (.A(_04636_),
    .X(clknet_0__04636_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04637_ (.A(_04637_),
    .X(clknet_0__04637_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04638_ (.A(_04638_),
    .X(clknet_0__04638_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04639_ (.A(_04639_),
    .X(clknet_0__04639_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04640_ (.A(_04640_),
    .X(clknet_0__04640_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04641_ (.A(_04641_),
    .X(clknet_0__04641_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04642_ (.A(_04642_),
    .X(clknet_0__04642_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04643_ (.A(_04643_),
    .X(clknet_0__04643_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04644_ (.A(_04644_),
    .X(clknet_0__04644_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04645_ (.A(_04645_),
    .X(clknet_0__04645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04646_ (.A(_04646_),
    .X(clknet_0__04646_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04647_ (.A(_04647_),
    .X(clknet_0__04647_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04648_ (.A(_04648_),
    .X(clknet_0__04648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04649_ (.A(_04649_),
    .X(clknet_0__04649_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04650_ (.A(_04650_),
    .X(clknet_0__04650_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04651_ (.A(_04651_),
    .X(clknet_0__04651_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04652_ (.A(_04652_),
    .X(clknet_0__04652_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04653_ (.A(_04653_),
    .X(clknet_0__04653_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04658_ (.A(_04658_),
    .X(clknet_0__04658_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04659_ (.A(_04659_),
    .X(clknet_0__04659_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04664_ (.A(_04664_),
    .X(clknet_0__04664_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04665_ (.A(_04665_),
    .X(clknet_0__04665_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04670_ (.A(_04670_),
    .X(clknet_0__04670_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04671_ (.A(_04671_),
    .X(clknet_0__04671_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04672_ (.A(_04672_),
    .X(clknet_0__04672_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04673_ (.A(_04673_),
    .X(clknet_0__04673_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04674_ (.A(_04674_),
    .X(clknet_0__04674_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04675_ (.A(_04675_),
    .X(clknet_0__04675_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04676_ (.A(_04676_),
    .X(clknet_0__04676_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04679_ (.A(_04679_),
    .X(clknet_0__04679_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04680_ (.A(_04680_),
    .X(clknet_0__04680_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04682_ (.A(_04682_),
    .X(clknet_0__04682_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04685_ (.A(_04685_),
    .X(clknet_0__04685_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0__04686_ (.A(_04686_),
    .X(clknet_0__04686_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_mclk (.A(net1692),
    .X(clknet_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock1 (.A(user_clock1),
    .X(clknet_0_user_clock1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_user_clock2 (.A(user_clock2),
    .X(clknet_0_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04347_ (.A(clknet_0__04347_),
    .X(clknet_1_0__leaf__04347_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04354_ (.A(clknet_0__04354_),
    .X(clknet_1_0__leaf__04354_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04355_ (.A(clknet_0__04355_),
    .X(clknet_1_0__leaf__04355_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04356_ (.A(clknet_0__04356_),
    .X(clknet_1_0__leaf__04356_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04357_ (.A(clknet_0__04357_),
    .X(clknet_1_0__leaf__04357_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04392_ (.A(clknet_0__04392_),
    .X(clknet_1_0__leaf__04392_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04393_ (.A(clknet_0__04393_),
    .X(clknet_1_0__leaf__04393_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04394_ (.A(clknet_0__04394_),
    .X(clknet_1_0__leaf__04394_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04395_ (.A(clknet_0__04395_),
    .X(clknet_1_0__leaf__04395_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04396_ (.A(clknet_0__04396_),
    .X(clknet_1_0__leaf__04396_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04397_ (.A(clknet_0__04397_),
    .X(clknet_1_0__leaf__04397_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04398_ (.A(clknet_0__04398_),
    .X(clknet_1_0__leaf__04398_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04399_ (.A(clknet_0__04399_),
    .X(clknet_1_0__leaf__04399_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04400_ (.A(clknet_0__04400_),
    .X(clknet_1_0__leaf__04400_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04401_ (.A(clknet_0__04401_),
    .X(clknet_1_0__leaf__04401_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04402_ (.A(clknet_0__04402_),
    .X(clknet_1_0__leaf__04402_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04403_ (.A(clknet_0__04403_),
    .X(clknet_1_0__leaf__04403_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04404_ (.A(clknet_0__04404_),
    .X(clknet_1_0__leaf__04404_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04405_ (.A(clknet_0__04405_),
    .X(clknet_1_0__leaf__04405_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04406_ (.A(clknet_0__04406_),
    .X(clknet_1_0__leaf__04406_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04407_ (.A(clknet_0__04407_),
    .X(clknet_1_0__leaf__04407_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04408_ (.A(clknet_0__04408_),
    .X(clknet_1_0__leaf__04408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04409_ (.A(clknet_0__04409_),
    .X(clknet_1_0__leaf__04409_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04410_ (.A(clknet_0__04410_),
    .X(clknet_1_0__leaf__04410_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04411_ (.A(clknet_0__04411_),
    .X(clknet_1_0__leaf__04411_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04412_ (.A(clknet_0__04412_),
    .X(clknet_1_0__leaf__04412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04413_ (.A(clknet_0__04413_),
    .X(clknet_1_0__leaf__04413_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04414_ (.A(clknet_0__04414_),
    .X(clknet_1_0__leaf__04414_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04415_ (.A(clknet_0__04415_),
    .X(clknet_1_0__leaf__04415_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04416_ (.A(clknet_0__04416_),
    .X(clknet_1_0__leaf__04416_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04417_ (.A(clknet_0__04417_),
    .X(clknet_1_0__leaf__04417_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04418_ (.A(clknet_0__04418_),
    .X(clknet_1_0__leaf__04418_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04419_ (.A(clknet_0__04419_),
    .X(clknet_1_0__leaf__04419_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04420_ (.A(clknet_0__04420_),
    .X(clknet_1_0__leaf__04420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04421_ (.A(clknet_0__04421_),
    .X(clknet_1_0__leaf__04421_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04422_ (.A(clknet_0__04422_),
    .X(clknet_1_0__leaf__04422_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04423_ (.A(clknet_0__04423_),
    .X(clknet_1_0__leaf__04423_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04424_ (.A(clknet_0__04424_),
    .X(clknet_1_0__leaf__04424_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04425_ (.A(clknet_0__04425_),
    .X(clknet_1_0__leaf__04425_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04426_ (.A(clknet_0__04426_),
    .X(clknet_1_0__leaf__04426_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04427_ (.A(clknet_0__04427_),
    .X(clknet_1_0__leaf__04427_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04428_ (.A(clknet_0__04428_),
    .X(clknet_1_0__leaf__04428_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04429_ (.A(clknet_0__04429_),
    .X(clknet_1_0__leaf__04429_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04430_ (.A(clknet_0__04430_),
    .X(clknet_1_0__leaf__04430_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04431_ (.A(clknet_0__04431_),
    .X(clknet_1_0__leaf__04431_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04432_ (.A(clknet_0__04432_),
    .X(clknet_1_0__leaf__04432_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04433_ (.A(clknet_0__04433_),
    .X(clknet_1_0__leaf__04433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04434_ (.A(clknet_0__04434_),
    .X(clknet_1_0__leaf__04434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04435_ (.A(clknet_0__04435_),
    .X(clknet_1_0__leaf__04435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04436_ (.A(clknet_0__04436_),
    .X(clknet_1_0__leaf__04436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04437_ (.A(clknet_0__04437_),
    .X(clknet_1_0__leaf__04437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04438_ (.A(clknet_0__04438_),
    .X(clknet_1_0__leaf__04438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04439_ (.A(clknet_0__04439_),
    .X(clknet_1_0__leaf__04439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04440_ (.A(clknet_0__04440_),
    .X(clknet_1_0__leaf__04440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04441_ (.A(clknet_0__04441_),
    .X(clknet_1_0__leaf__04441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04442_ (.A(clknet_0__04442_),
    .X(clknet_1_0__leaf__04442_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04443_ (.A(clknet_0__04443_),
    .X(clknet_1_0__leaf__04443_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04444_ (.A(clknet_0__04444_),
    .X(clknet_1_0__leaf__04444_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04445_ (.A(clknet_0__04445_),
    .X(clknet_1_0__leaf__04445_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04446_ (.A(clknet_0__04446_),
    .X(clknet_1_0__leaf__04446_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04447_ (.A(clknet_0__04447_),
    .X(clknet_1_0__leaf__04447_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04448_ (.A(clknet_0__04448_),
    .X(clknet_1_0__leaf__04448_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04449_ (.A(clknet_0__04449_),
    .X(clknet_1_0__leaf__04449_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04450_ (.A(clknet_0__04450_),
    .X(clknet_1_0__leaf__04450_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04451_ (.A(clknet_0__04451_),
    .X(clknet_1_0__leaf__04451_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04452_ (.A(clknet_0__04452_),
    .X(clknet_1_0__leaf__04452_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04453_ (.A(clknet_0__04453_),
    .X(clknet_1_0__leaf__04453_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04454_ (.A(clknet_0__04454_),
    .X(clknet_1_0__leaf__04454_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04455_ (.A(clknet_0__04455_),
    .X(clknet_1_0__leaf__04455_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04456_ (.A(clknet_0__04456_),
    .X(clknet_1_0__leaf__04456_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04457_ (.A(clknet_0__04457_),
    .X(clknet_1_0__leaf__04457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04458_ (.A(clknet_0__04458_),
    .X(clknet_1_0__leaf__04458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04459_ (.A(clknet_0__04459_),
    .X(clknet_1_0__leaf__04459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04460_ (.A(clknet_0__04460_),
    .X(clknet_1_0__leaf__04460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04461_ (.A(clknet_0__04461_),
    .X(clknet_1_0__leaf__04461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04463_ (.A(clknet_0__04463_),
    .X(clknet_1_0__leaf__04463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04464_ (.A(clknet_0__04464_),
    .X(clknet_1_0__leaf__04464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04465_ (.A(clknet_0__04465_),
    .X(clknet_1_0__leaf__04465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04466_ (.A(clknet_0__04466_),
    .X(clknet_1_0__leaf__04466_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04467_ (.A(clknet_0__04467_),
    .X(clknet_1_0__leaf__04467_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04468_ (.A(clknet_0__04468_),
    .X(clknet_1_0__leaf__04468_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04469_ (.A(clknet_0__04469_),
    .X(clknet_1_0__leaf__04469_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04470_ (.A(clknet_0__04470_),
    .X(clknet_1_0__leaf__04470_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04471_ (.A(clknet_0__04471_),
    .X(clknet_1_0__leaf__04471_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04472_ (.A(clknet_0__04472_),
    .X(clknet_1_0__leaf__04472_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04473_ (.A(clknet_0__04473_),
    .X(clknet_1_0__leaf__04473_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04474_ (.A(clknet_0__04474_),
    .X(clknet_1_0__leaf__04474_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04475_ (.A(clknet_0__04475_),
    .X(clknet_1_0__leaf__04475_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04476_ (.A(clknet_0__04476_),
    .X(clknet_1_0__leaf__04476_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04477_ (.A(clknet_0__04477_),
    .X(clknet_1_0__leaf__04477_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04478_ (.A(clknet_0__04478_),
    .X(clknet_1_0__leaf__04478_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04479_ (.A(clknet_0__04479_),
    .X(clknet_1_0__leaf__04479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04480_ (.A(clknet_0__04480_),
    .X(clknet_1_0__leaf__04480_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04481_ (.A(clknet_0__04481_),
    .X(clknet_1_0__leaf__04481_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04482_ (.A(clknet_0__04482_),
    .X(clknet_1_0__leaf__04482_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04483_ (.A(clknet_0__04483_),
    .X(clknet_1_0__leaf__04483_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04484_ (.A(clknet_0__04484_),
    .X(clknet_1_0__leaf__04484_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04485_ (.A(clknet_0__04485_),
    .X(clknet_1_0__leaf__04485_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04486_ (.A(clknet_0__04486_),
    .X(clknet_1_0__leaf__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04487_ (.A(clknet_0__04487_),
    .X(clknet_1_0__leaf__04487_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04488_ (.A(clknet_0__04488_),
    .X(clknet_1_0__leaf__04488_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04489_ (.A(clknet_0__04489_),
    .X(clknet_1_0__leaf__04489_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04490_ (.A(clknet_0__04490_),
    .X(clknet_1_0__leaf__04490_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04491_ (.A(clknet_0__04491_),
    .X(clknet_1_0__leaf__04491_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04492_ (.A(clknet_0__04492_),
    .X(clknet_1_0__leaf__04492_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04494_ (.A(clknet_0__04494_),
    .X(clknet_1_0__leaf__04494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04495_ (.A(clknet_0__04495_),
    .X(clknet_1_0__leaf__04495_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04496_ (.A(clknet_0__04496_),
    .X(clknet_1_0__leaf__04496_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04497_ (.A(clknet_0__04497_),
    .X(clknet_1_0__leaf__04497_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04498_ (.A(clknet_0__04498_),
    .X(clknet_1_0__leaf__04498_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04499_ (.A(clknet_0__04499_),
    .X(clknet_1_0__leaf__04499_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04500_ (.A(clknet_0__04500_),
    .X(clknet_1_0__leaf__04500_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04501_ (.A(clknet_0__04501_),
    .X(clknet_1_0__leaf__04501_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04502_ (.A(clknet_0__04502_),
    .X(clknet_1_0__leaf__04502_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04503_ (.A(clknet_0__04503_),
    .X(clknet_1_0__leaf__04503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04504_ (.A(clknet_0__04504_),
    .X(clknet_1_0__leaf__04504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04505_ (.A(clknet_0__04505_),
    .X(clknet_1_0__leaf__04505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04538_ (.A(clknet_0__04538_),
    .X(clknet_1_0__leaf__04538_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04539_ (.A(clknet_0__04539_),
    .X(clknet_1_0__leaf__04539_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04540_ (.A(clknet_0__04540_),
    .X(clknet_1_0__leaf__04540_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04541_ (.A(clknet_0__04541_),
    .X(clknet_1_0__leaf__04541_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04542_ (.A(clknet_0__04542_),
    .X(clknet_1_0__leaf__04542_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04543_ (.A(clknet_0__04543_),
    .X(clknet_1_0__leaf__04543_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04544_ (.A(clknet_0__04544_),
    .X(clknet_1_0__leaf__04544_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04545_ (.A(clknet_0__04545_),
    .X(clknet_1_0__leaf__04545_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04546_ (.A(clknet_0__04546_),
    .X(clknet_1_0__leaf__04546_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04547_ (.A(clknet_0__04547_),
    .X(clknet_1_0__leaf__04547_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04548_ (.A(clknet_0__04548_),
    .X(clknet_1_0__leaf__04548_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04549_ (.A(clknet_0__04549_),
    .X(clknet_1_0__leaf__04549_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04550_ (.A(clknet_0__04550_),
    .X(clknet_1_0__leaf__04550_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04551_ (.A(clknet_0__04551_),
    .X(clknet_1_0__leaf__04551_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04552_ (.A(clknet_0__04552_),
    .X(clknet_1_0__leaf__04552_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04562_ (.A(clknet_0__04562_),
    .X(clknet_1_0__leaf__04562_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04565_ (.A(clknet_0__04565_),
    .X(clknet_1_0__leaf__04565_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04566_ (.A(clknet_0__04566_),
    .X(clknet_1_0__leaf__04566_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04568_ (.A(clknet_0__04568_),
    .X(clknet_1_0__leaf__04568_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04569_ (.A(clknet_0__04569_),
    .X(clknet_1_0__leaf__04569_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04570_ (.A(clknet_0__04570_),
    .X(clknet_1_0__leaf__04570_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04571_ (.A(clknet_0__04571_),
    .X(clknet_1_0__leaf__04571_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04572_ (.A(clknet_0__04572_),
    .X(clknet_1_0__leaf__04572_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04573_ (.A(clknet_0__04573_),
    .X(clknet_1_0__leaf__04573_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04574_ (.A(clknet_0__04574_),
    .X(clknet_1_0__leaf__04574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04575_ (.A(clknet_0__04575_),
    .X(clknet_1_0__leaf__04575_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04576_ (.A(clknet_0__04576_),
    .X(clknet_1_0__leaf__04576_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04577_ (.A(clknet_0__04577_),
    .X(clknet_1_0__leaf__04577_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04578_ (.A(clknet_0__04578_),
    .X(clknet_1_0__leaf__04578_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04579_ (.A(clknet_0__04579_),
    .X(clknet_1_0__leaf__04579_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04580_ (.A(clknet_0__04580_),
    .X(clknet_1_0__leaf__04580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04581_ (.A(clknet_0__04581_),
    .X(clknet_1_0__leaf__04581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04582_ (.A(clknet_0__04582_),
    .X(clknet_1_0__leaf__04582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04583_ (.A(clknet_0__04583_),
    .X(clknet_1_0__leaf__04583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04584_ (.A(clknet_0__04584_),
    .X(clknet_1_0__leaf__04584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04587_ (.A(clknet_0__04587_),
    .X(clknet_1_0__leaf__04587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04588_ (.A(clknet_0__04588_),
    .X(clknet_1_0__leaf__04588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04590_ (.A(clknet_0__04590_),
    .X(clknet_1_0__leaf__04590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04591_ (.A(clknet_0__04591_),
    .X(clknet_1_0__leaf__04591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04592_ (.A(clknet_0__04592_),
    .X(clknet_1_0__leaf__04592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04593_ (.A(clknet_0__04593_),
    .X(clknet_1_0__leaf__04593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04594_ (.A(clknet_0__04594_),
    .X(clknet_1_0__leaf__04594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04595_ (.A(clknet_0__04595_),
    .X(clknet_1_0__leaf__04595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04596_ (.A(clknet_0__04596_),
    .X(clknet_1_0__leaf__04596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04597_ (.A(clknet_0__04597_),
    .X(clknet_1_0__leaf__04597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04598_ (.A(clknet_0__04598_),
    .X(clknet_1_0__leaf__04598_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04599_ (.A(clknet_0__04599_),
    .X(clknet_1_0__leaf__04599_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04600_ (.A(clknet_0__04600_),
    .X(clknet_1_0__leaf__04600_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04601_ (.A(clknet_0__04601_),
    .X(clknet_1_0__leaf__04601_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04602_ (.A(clknet_0__04602_),
    .X(clknet_1_0__leaf__04602_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04603_ (.A(clknet_0__04603_),
    .X(clknet_1_0__leaf__04603_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04604_ (.A(clknet_0__04604_),
    .X(clknet_1_0__leaf__04604_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04605_ (.A(clknet_0__04605_),
    .X(clknet_1_0__leaf__04605_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04606_ (.A(clknet_0__04606_),
    .X(clknet_1_0__leaf__04606_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04609_ (.A(clknet_0__04609_),
    .X(clknet_1_0__leaf__04609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04610_ (.A(clknet_0__04610_),
    .X(clknet_1_0__leaf__04610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04612_ (.A(clknet_0__04612_),
    .X(clknet_1_0__leaf__04612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04613_ (.A(clknet_0__04613_),
    .X(clknet_1_0__leaf__04613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04614_ (.A(clknet_0__04614_),
    .X(clknet_1_0__leaf__04614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04615_ (.A(clknet_0__04615_),
    .X(clknet_1_0__leaf__04615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04616_ (.A(clknet_0__04616_),
    .X(clknet_1_0__leaf__04616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04617_ (.A(clknet_0__04617_),
    .X(clknet_1_0__leaf__04617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04618_ (.A(clknet_0__04618_),
    .X(clknet_1_0__leaf__04618_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04619_ (.A(clknet_0__04619_),
    .X(clknet_1_0__leaf__04619_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04620_ (.A(clknet_0__04620_),
    .X(clknet_1_0__leaf__04620_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04621_ (.A(clknet_0__04621_),
    .X(clknet_1_0__leaf__04621_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04622_ (.A(clknet_0__04622_),
    .X(clknet_1_0__leaf__04622_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04623_ (.A(clknet_0__04623_),
    .X(clknet_1_0__leaf__04623_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04624_ (.A(clknet_0__04624_),
    .X(clknet_1_0__leaf__04624_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04625_ (.A(clknet_0__04625_),
    .X(clknet_1_0__leaf__04625_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04626_ (.A(clknet_0__04626_),
    .X(clknet_1_0__leaf__04626_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04627_ (.A(clknet_0__04627_),
    .X(clknet_1_0__leaf__04627_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04628_ (.A(clknet_0__04628_),
    .X(clknet_1_0__leaf__04628_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04629_ (.A(clknet_0__04629_),
    .X(clknet_1_0__leaf__04629_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04630_ (.A(clknet_0__04630_),
    .X(clknet_1_0__leaf__04630_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04631_ (.A(clknet_0__04631_),
    .X(clknet_1_0__leaf__04631_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04632_ (.A(clknet_0__04632_),
    .X(clknet_1_0__leaf__04632_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04634_ (.A(clknet_0__04634_),
    .X(clknet_1_0__leaf__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04635_ (.A(clknet_0__04635_),
    .X(clknet_1_0__leaf__04635_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04636_ (.A(clknet_0__04636_),
    .X(clknet_1_0__leaf__04636_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04637_ (.A(clknet_0__04637_),
    .X(clknet_1_0__leaf__04637_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04638_ (.A(clknet_0__04638_),
    .X(clknet_1_0__leaf__04638_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04639_ (.A(clknet_0__04639_),
    .X(clknet_1_0__leaf__04639_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04640_ (.A(clknet_0__04640_),
    .X(clknet_1_0__leaf__04640_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04641_ (.A(clknet_0__04641_),
    .X(clknet_1_0__leaf__04641_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04642_ (.A(clknet_0__04642_),
    .X(clknet_1_0__leaf__04642_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04643_ (.A(clknet_0__04643_),
    .X(clknet_1_0__leaf__04643_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04644_ (.A(clknet_0__04644_),
    .X(clknet_1_0__leaf__04644_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04645_ (.A(clknet_0__04645_),
    .X(clknet_1_0__leaf__04645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04646_ (.A(clknet_0__04646_),
    .X(clknet_1_0__leaf__04646_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04647_ (.A(clknet_0__04647_),
    .X(clknet_1_0__leaf__04647_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04648_ (.A(clknet_0__04648_),
    .X(clknet_1_0__leaf__04648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04649_ (.A(clknet_0__04649_),
    .X(clknet_1_0__leaf__04649_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04650_ (.A(clknet_0__04650_),
    .X(clknet_1_0__leaf__04650_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04651_ (.A(clknet_0__04651_),
    .X(clknet_1_0__leaf__04651_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04652_ (.A(clknet_0__04652_),
    .X(clknet_1_0__leaf__04652_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04658_ (.A(clknet_0__04658_),
    .X(clknet_1_0__leaf__04658_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04659_ (.A(clknet_0__04659_),
    .X(clknet_1_0__leaf__04659_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04664_ (.A(clknet_0__04664_),
    .X(clknet_1_0__leaf__04664_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04665_ (.A(clknet_0__04665_),
    .X(clknet_1_0__leaf__04665_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04670_ (.A(clknet_0__04670_),
    .X(clknet_1_0__leaf__04670_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04671_ (.A(clknet_0__04671_),
    .X(clknet_1_0__leaf__04671_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04672_ (.A(clknet_0__04672_),
    .X(clknet_1_0__leaf__04672_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04673_ (.A(clknet_0__04673_),
    .X(clknet_1_0__leaf__04673_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04674_ (.A(clknet_0__04674_),
    .X(clknet_1_0__leaf__04674_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04675_ (.A(clknet_0__04675_),
    .X(clknet_1_0__leaf__04675_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04676_ (.A(clknet_0__04676_),
    .X(clknet_1_0__leaf__04676_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04679_ (.A(clknet_0__04679_),
    .X(clknet_1_0__leaf__04679_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04680_ (.A(clknet_0__04680_),
    .X(clknet_1_0__leaf__04680_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04682_ (.A(clknet_0__04682_),
    .X(clknet_1_0__leaf__04682_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04685_ (.A(clknet_0__04685_),
    .X(clknet_1_0__leaf__04685_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f__04686_ (.A(clknet_0__04686_),
    .X(clknet_1_0__leaf__04686_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_user_clock1 (.A(clknet_0_user_clock1),
    .X(clknet_1_0__leaf_user_clock1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_0__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04347_ (.A(clknet_0__04347_),
    .X(clknet_1_1__leaf__04347_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04354_ (.A(clknet_0__04354_),
    .X(clknet_1_1__leaf__04354_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04355_ (.A(clknet_0__04355_),
    .X(clknet_1_1__leaf__04355_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04356_ (.A(clknet_0__04356_),
    .X(clknet_1_1__leaf__04356_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04357_ (.A(clknet_0__04357_),
    .X(clknet_1_1__leaf__04357_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04392_ (.A(clknet_0__04392_),
    .X(clknet_1_1__leaf__04392_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04393_ (.A(clknet_0__04393_),
    .X(clknet_1_1__leaf__04393_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04394_ (.A(clknet_0__04394_),
    .X(clknet_1_1__leaf__04394_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04395_ (.A(clknet_0__04395_),
    .X(clknet_1_1__leaf__04395_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04396_ (.A(clknet_0__04396_),
    .X(clknet_1_1__leaf__04396_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04397_ (.A(clknet_0__04397_),
    .X(clknet_1_1__leaf__04397_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04398_ (.A(clknet_0__04398_),
    .X(clknet_1_1__leaf__04398_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04399_ (.A(clknet_0__04399_),
    .X(clknet_1_1__leaf__04399_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04400_ (.A(clknet_0__04400_),
    .X(clknet_1_1__leaf__04400_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04401_ (.A(clknet_0__04401_),
    .X(clknet_1_1__leaf__04401_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04402_ (.A(clknet_0__04402_),
    .X(clknet_1_1__leaf__04402_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04403_ (.A(clknet_0__04403_),
    .X(clknet_1_1__leaf__04403_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04404_ (.A(clknet_0__04404_),
    .X(clknet_1_1__leaf__04404_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04405_ (.A(clknet_0__04405_),
    .X(clknet_1_1__leaf__04405_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04406_ (.A(clknet_0__04406_),
    .X(clknet_1_1__leaf__04406_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04407_ (.A(clknet_0__04407_),
    .X(clknet_1_1__leaf__04407_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04408_ (.A(clknet_0__04408_),
    .X(clknet_1_1__leaf__04408_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04409_ (.A(clknet_0__04409_),
    .X(clknet_1_1__leaf__04409_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04410_ (.A(clknet_0__04410_),
    .X(clknet_1_1__leaf__04410_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04411_ (.A(clknet_0__04411_),
    .X(clknet_1_1__leaf__04411_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04412_ (.A(clknet_0__04412_),
    .X(clknet_1_1__leaf__04412_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04413_ (.A(clknet_0__04413_),
    .X(clknet_1_1__leaf__04413_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04414_ (.A(clknet_0__04414_),
    .X(clknet_1_1__leaf__04414_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04415_ (.A(clknet_0__04415_),
    .X(clknet_1_1__leaf__04415_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04416_ (.A(clknet_0__04416_),
    .X(clknet_1_1__leaf__04416_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04417_ (.A(clknet_0__04417_),
    .X(clknet_1_1__leaf__04417_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04418_ (.A(clknet_0__04418_),
    .X(clknet_1_1__leaf__04418_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04419_ (.A(clknet_0__04419_),
    .X(clknet_1_1__leaf__04419_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04420_ (.A(clknet_0__04420_),
    .X(clknet_1_1__leaf__04420_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04421_ (.A(clknet_0__04421_),
    .X(clknet_1_1__leaf__04421_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04422_ (.A(clknet_0__04422_),
    .X(clknet_1_1__leaf__04422_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04423_ (.A(clknet_0__04423_),
    .X(clknet_1_1__leaf__04423_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04424_ (.A(clknet_0__04424_),
    .X(clknet_1_1__leaf__04424_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04425_ (.A(clknet_0__04425_),
    .X(clknet_1_1__leaf__04425_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04426_ (.A(clknet_0__04426_),
    .X(clknet_1_1__leaf__04426_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04427_ (.A(clknet_0__04427_),
    .X(clknet_1_1__leaf__04427_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04428_ (.A(clknet_0__04428_),
    .X(clknet_1_1__leaf__04428_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04429_ (.A(clknet_0__04429_),
    .X(clknet_1_1__leaf__04429_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04430_ (.A(clknet_0__04430_),
    .X(clknet_1_1__leaf__04430_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04431_ (.A(clknet_0__04431_),
    .X(clknet_1_1__leaf__04431_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04432_ (.A(clknet_0__04432_),
    .X(clknet_1_1__leaf__04432_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04433_ (.A(clknet_0__04433_),
    .X(clknet_1_1__leaf__04433_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04434_ (.A(clknet_0__04434_),
    .X(clknet_1_1__leaf__04434_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04435_ (.A(clknet_0__04435_),
    .X(clknet_1_1__leaf__04435_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04436_ (.A(clknet_0__04436_),
    .X(clknet_1_1__leaf__04436_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04437_ (.A(clknet_0__04437_),
    .X(clknet_1_1__leaf__04437_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04438_ (.A(clknet_0__04438_),
    .X(clknet_1_1__leaf__04438_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04439_ (.A(clknet_0__04439_),
    .X(clknet_1_1__leaf__04439_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04440_ (.A(clknet_0__04440_),
    .X(clknet_1_1__leaf__04440_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04441_ (.A(clknet_0__04441_),
    .X(clknet_1_1__leaf__04441_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04442_ (.A(clknet_0__04442_),
    .X(clknet_1_1__leaf__04442_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04443_ (.A(clknet_0__04443_),
    .X(clknet_1_1__leaf__04443_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04444_ (.A(clknet_0__04444_),
    .X(clknet_1_1__leaf__04444_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04445_ (.A(clknet_0__04445_),
    .X(clknet_1_1__leaf__04445_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04446_ (.A(clknet_0__04446_),
    .X(clknet_1_1__leaf__04446_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04447_ (.A(clknet_0__04447_),
    .X(clknet_1_1__leaf__04447_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04448_ (.A(clknet_0__04448_),
    .X(clknet_1_1__leaf__04448_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04449_ (.A(clknet_0__04449_),
    .X(clknet_1_1__leaf__04449_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04450_ (.A(clknet_0__04450_),
    .X(clknet_1_1__leaf__04450_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04451_ (.A(clknet_0__04451_),
    .X(clknet_1_1__leaf__04451_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04452_ (.A(clknet_0__04452_),
    .X(clknet_1_1__leaf__04452_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04453_ (.A(clknet_0__04453_),
    .X(clknet_1_1__leaf__04453_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04454_ (.A(clknet_0__04454_),
    .X(clknet_1_1__leaf__04454_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04455_ (.A(clknet_0__04455_),
    .X(clknet_1_1__leaf__04455_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04456_ (.A(clknet_0__04456_),
    .X(clknet_1_1__leaf__04456_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04457_ (.A(clknet_0__04457_),
    .X(clknet_1_1__leaf__04457_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04458_ (.A(clknet_0__04458_),
    .X(clknet_1_1__leaf__04458_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04459_ (.A(clknet_0__04459_),
    .X(clknet_1_1__leaf__04459_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04460_ (.A(clknet_0__04460_),
    .X(clknet_1_1__leaf__04460_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04461_ (.A(clknet_0__04461_),
    .X(clknet_1_1__leaf__04461_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04463_ (.A(clknet_0__04463_),
    .X(clknet_1_1__leaf__04463_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04464_ (.A(clknet_0__04464_),
    .X(clknet_1_1__leaf__04464_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04465_ (.A(clknet_0__04465_),
    .X(clknet_1_1__leaf__04465_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04466_ (.A(clknet_0__04466_),
    .X(clknet_1_1__leaf__04466_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04467_ (.A(clknet_0__04467_),
    .X(clknet_1_1__leaf__04467_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04468_ (.A(clknet_0__04468_),
    .X(clknet_1_1__leaf__04468_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04469_ (.A(clknet_0__04469_),
    .X(clknet_1_1__leaf__04469_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04470_ (.A(clknet_0__04470_),
    .X(clknet_1_1__leaf__04470_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04471_ (.A(clknet_0__04471_),
    .X(clknet_1_1__leaf__04471_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04472_ (.A(clknet_0__04472_),
    .X(clknet_1_1__leaf__04472_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04473_ (.A(clknet_0__04473_),
    .X(clknet_1_1__leaf__04473_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04474_ (.A(clknet_0__04474_),
    .X(clknet_1_1__leaf__04474_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04475_ (.A(clknet_0__04475_),
    .X(clknet_1_1__leaf__04475_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04476_ (.A(clknet_0__04476_),
    .X(clknet_1_1__leaf__04476_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04477_ (.A(clknet_0__04477_),
    .X(clknet_1_1__leaf__04477_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04478_ (.A(clknet_0__04478_),
    .X(clknet_1_1__leaf__04478_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04479_ (.A(clknet_0__04479_),
    .X(clknet_1_1__leaf__04479_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04480_ (.A(clknet_0__04480_),
    .X(clknet_1_1__leaf__04480_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04481_ (.A(clknet_0__04481_),
    .X(clknet_1_1__leaf__04481_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04482_ (.A(clknet_0__04482_),
    .X(clknet_1_1__leaf__04482_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04483_ (.A(clknet_0__04483_),
    .X(clknet_1_1__leaf__04483_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04484_ (.A(clknet_0__04484_),
    .X(clknet_1_1__leaf__04484_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04485_ (.A(clknet_0__04485_),
    .X(clknet_1_1__leaf__04485_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04486_ (.A(clknet_0__04486_),
    .X(clknet_1_1__leaf__04486_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04487_ (.A(clknet_0__04487_),
    .X(clknet_1_1__leaf__04487_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04488_ (.A(clknet_0__04488_),
    .X(clknet_1_1__leaf__04488_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04489_ (.A(clknet_0__04489_),
    .X(clknet_1_1__leaf__04489_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04490_ (.A(clknet_0__04490_),
    .X(clknet_1_1__leaf__04490_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04491_ (.A(clknet_0__04491_),
    .X(clknet_1_1__leaf__04491_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04492_ (.A(clknet_0__04492_),
    .X(clknet_1_1__leaf__04492_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04494_ (.A(clknet_0__04494_),
    .X(clknet_1_1__leaf__04494_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04495_ (.A(clknet_0__04495_),
    .X(clknet_1_1__leaf__04495_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04496_ (.A(clknet_0__04496_),
    .X(clknet_1_1__leaf__04496_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04497_ (.A(clknet_0__04497_),
    .X(clknet_1_1__leaf__04497_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04498_ (.A(clknet_0__04498_),
    .X(clknet_1_1__leaf__04498_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04499_ (.A(clknet_0__04499_),
    .X(clknet_1_1__leaf__04499_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04500_ (.A(clknet_0__04500_),
    .X(clknet_1_1__leaf__04500_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04501_ (.A(clknet_0__04501_),
    .X(clknet_1_1__leaf__04501_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04502_ (.A(clknet_0__04502_),
    .X(clknet_1_1__leaf__04502_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04503_ (.A(clknet_0__04503_),
    .X(clknet_1_1__leaf__04503_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04504_ (.A(clknet_0__04504_),
    .X(clknet_1_1__leaf__04504_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04505_ (.A(clknet_0__04505_),
    .X(clknet_1_1__leaf__04505_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04538_ (.A(clknet_0__04538_),
    .X(clknet_1_1__leaf__04538_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04539_ (.A(clknet_0__04539_),
    .X(clknet_1_1__leaf__04539_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04540_ (.A(clknet_0__04540_),
    .X(clknet_1_1__leaf__04540_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04541_ (.A(clknet_0__04541_),
    .X(clknet_1_1__leaf__04541_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04542_ (.A(clknet_0__04542_),
    .X(clknet_1_1__leaf__04542_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04543_ (.A(clknet_0__04543_),
    .X(clknet_1_1__leaf__04543_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04544_ (.A(clknet_0__04544_),
    .X(clknet_1_1__leaf__04544_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04545_ (.A(clknet_0__04545_),
    .X(clknet_1_1__leaf__04545_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04546_ (.A(clknet_0__04546_),
    .X(clknet_1_1__leaf__04546_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04547_ (.A(clknet_0__04547_),
    .X(clknet_1_1__leaf__04547_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04548_ (.A(clknet_0__04548_),
    .X(clknet_1_1__leaf__04548_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04549_ (.A(clknet_0__04549_),
    .X(clknet_1_1__leaf__04549_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04550_ (.A(clknet_0__04550_),
    .X(clknet_1_1__leaf__04550_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04551_ (.A(clknet_0__04551_),
    .X(clknet_1_1__leaf__04551_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04552_ (.A(clknet_0__04552_),
    .X(clknet_1_1__leaf__04552_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04562_ (.A(clknet_0__04562_),
    .X(clknet_1_1__leaf__04562_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04565_ (.A(clknet_0__04565_),
    .X(clknet_1_1__leaf__04565_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04566_ (.A(clknet_0__04566_),
    .X(clknet_1_1__leaf__04566_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04568_ (.A(clknet_0__04568_),
    .X(clknet_1_1__leaf__04568_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04569_ (.A(clknet_0__04569_),
    .X(clknet_1_1__leaf__04569_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04570_ (.A(clknet_0__04570_),
    .X(clknet_1_1__leaf__04570_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04571_ (.A(clknet_0__04571_),
    .X(clknet_1_1__leaf__04571_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04572_ (.A(clknet_0__04572_),
    .X(clknet_1_1__leaf__04572_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04573_ (.A(clknet_0__04573_),
    .X(clknet_1_1__leaf__04573_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04574_ (.A(clknet_0__04574_),
    .X(clknet_1_1__leaf__04574_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04575_ (.A(clknet_0__04575_),
    .X(clknet_1_1__leaf__04575_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04576_ (.A(clknet_0__04576_),
    .X(clknet_1_1__leaf__04576_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04577_ (.A(clknet_0__04577_),
    .X(clknet_1_1__leaf__04577_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04578_ (.A(clknet_0__04578_),
    .X(clknet_1_1__leaf__04578_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04579_ (.A(clknet_0__04579_),
    .X(clknet_1_1__leaf__04579_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04580_ (.A(clknet_0__04580_),
    .X(clknet_1_1__leaf__04580_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04581_ (.A(clknet_0__04581_),
    .X(clknet_1_1__leaf__04581_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04582_ (.A(clknet_0__04582_),
    .X(clknet_1_1__leaf__04582_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04583_ (.A(clknet_0__04583_),
    .X(clknet_1_1__leaf__04583_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04584_ (.A(clknet_0__04584_),
    .X(clknet_1_1__leaf__04584_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04587_ (.A(clknet_0__04587_),
    .X(clknet_1_1__leaf__04587_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04588_ (.A(clknet_0__04588_),
    .X(clknet_1_1__leaf__04588_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04590_ (.A(clknet_0__04590_),
    .X(clknet_1_1__leaf__04590_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04591_ (.A(clknet_0__04591_),
    .X(clknet_1_1__leaf__04591_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04592_ (.A(clknet_0__04592_),
    .X(clknet_1_1__leaf__04592_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04593_ (.A(clknet_0__04593_),
    .X(clknet_1_1__leaf__04593_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04594_ (.A(clknet_0__04594_),
    .X(clknet_1_1__leaf__04594_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04595_ (.A(clknet_0__04595_),
    .X(clknet_1_1__leaf__04595_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04596_ (.A(clknet_0__04596_),
    .X(clknet_1_1__leaf__04596_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04597_ (.A(clknet_0__04597_),
    .X(clknet_1_1__leaf__04597_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04598_ (.A(clknet_0__04598_),
    .X(clknet_1_1__leaf__04598_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04599_ (.A(clknet_0__04599_),
    .X(clknet_1_1__leaf__04599_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04600_ (.A(clknet_0__04600_),
    .X(clknet_1_1__leaf__04600_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04601_ (.A(clknet_0__04601_),
    .X(clknet_1_1__leaf__04601_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04602_ (.A(clknet_0__04602_),
    .X(clknet_1_1__leaf__04602_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04603_ (.A(clknet_0__04603_),
    .X(clknet_1_1__leaf__04603_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04604_ (.A(clknet_0__04604_),
    .X(clknet_1_1__leaf__04604_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04605_ (.A(clknet_0__04605_),
    .X(clknet_1_1__leaf__04605_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04606_ (.A(clknet_0__04606_),
    .X(clknet_1_1__leaf__04606_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04609_ (.A(clknet_0__04609_),
    .X(clknet_1_1__leaf__04609_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04610_ (.A(clknet_0__04610_),
    .X(clknet_1_1__leaf__04610_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04612_ (.A(clknet_0__04612_),
    .X(clknet_1_1__leaf__04612_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04613_ (.A(clknet_0__04613_),
    .X(clknet_1_1__leaf__04613_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04614_ (.A(clknet_0__04614_),
    .X(clknet_1_1__leaf__04614_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04615_ (.A(clknet_0__04615_),
    .X(clknet_1_1__leaf__04615_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04616_ (.A(clknet_0__04616_),
    .X(clknet_1_1__leaf__04616_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04617_ (.A(clknet_0__04617_),
    .X(clknet_1_1__leaf__04617_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04618_ (.A(clknet_0__04618_),
    .X(clknet_1_1__leaf__04618_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04619_ (.A(clknet_0__04619_),
    .X(clknet_1_1__leaf__04619_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04620_ (.A(clknet_0__04620_),
    .X(clknet_1_1__leaf__04620_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04621_ (.A(clknet_0__04621_),
    .X(clknet_1_1__leaf__04621_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04622_ (.A(clknet_0__04622_),
    .X(clknet_1_1__leaf__04622_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04623_ (.A(clknet_0__04623_),
    .X(clknet_1_1__leaf__04623_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04624_ (.A(clknet_0__04624_),
    .X(clknet_1_1__leaf__04624_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04625_ (.A(clknet_0__04625_),
    .X(clknet_1_1__leaf__04625_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04626_ (.A(clknet_0__04626_),
    .X(clknet_1_1__leaf__04626_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04627_ (.A(clknet_0__04627_),
    .X(clknet_1_1__leaf__04627_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04628_ (.A(clknet_0__04628_),
    .X(clknet_1_1__leaf__04628_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04629_ (.A(clknet_0__04629_),
    .X(clknet_1_1__leaf__04629_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04630_ (.A(clknet_0__04630_),
    .X(clknet_1_1__leaf__04630_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04631_ (.A(clknet_0__04631_),
    .X(clknet_1_1__leaf__04631_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04632_ (.A(clknet_0__04632_),
    .X(clknet_1_1__leaf__04632_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04634_ (.A(clknet_0__04634_),
    .X(clknet_1_1__leaf__04634_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04635_ (.A(clknet_0__04635_),
    .X(clknet_1_1__leaf__04635_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04636_ (.A(clknet_0__04636_),
    .X(clknet_1_1__leaf__04636_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04637_ (.A(clknet_0__04637_),
    .X(clknet_1_1__leaf__04637_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04638_ (.A(clknet_0__04638_),
    .X(clknet_1_1__leaf__04638_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04639_ (.A(clknet_0__04639_),
    .X(clknet_1_1__leaf__04639_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04640_ (.A(clknet_0__04640_),
    .X(clknet_1_1__leaf__04640_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04641_ (.A(clknet_0__04641_),
    .X(clknet_1_1__leaf__04641_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04642_ (.A(clknet_0__04642_),
    .X(clknet_1_1__leaf__04642_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04643_ (.A(clknet_0__04643_),
    .X(clknet_1_1__leaf__04643_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04644_ (.A(clknet_0__04644_),
    .X(clknet_1_1__leaf__04644_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04645_ (.A(clknet_0__04645_),
    .X(clknet_1_1__leaf__04645_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04646_ (.A(clknet_0__04646_),
    .X(clknet_1_1__leaf__04646_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04647_ (.A(clknet_0__04647_),
    .X(clknet_1_1__leaf__04647_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04648_ (.A(clknet_0__04648_),
    .X(clknet_1_1__leaf__04648_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04649_ (.A(clknet_0__04649_),
    .X(clknet_1_1__leaf__04649_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04650_ (.A(clknet_0__04650_),
    .X(clknet_1_1__leaf__04650_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04651_ (.A(clknet_0__04651_),
    .X(clknet_1_1__leaf__04651_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04652_ (.A(clknet_0__04652_),
    .X(clknet_1_1__leaf__04652_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04658_ (.A(clknet_0__04658_),
    .X(clknet_1_1__leaf__04658_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04659_ (.A(clknet_0__04659_),
    .X(clknet_1_1__leaf__04659_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04664_ (.A(clknet_0__04664_),
    .X(clknet_1_1__leaf__04664_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04665_ (.A(clknet_0__04665_),
    .X(clknet_1_1__leaf__04665_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04670_ (.A(clknet_0__04670_),
    .X(clknet_1_1__leaf__04670_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04671_ (.A(clknet_0__04671_),
    .X(clknet_1_1__leaf__04671_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04672_ (.A(clknet_0__04672_),
    .X(clknet_1_1__leaf__04672_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04673_ (.A(clknet_0__04673_),
    .X(clknet_1_1__leaf__04673_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04674_ (.A(clknet_0__04674_),
    .X(clknet_1_1__leaf__04674_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04675_ (.A(clknet_0__04675_),
    .X(clknet_1_1__leaf__04675_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04676_ (.A(clknet_0__04676_),
    .X(clknet_1_1__leaf__04676_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04679_ (.A(clknet_0__04679_),
    .X(clknet_1_1__leaf__04679_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04680_ (.A(clknet_0__04680_),
    .X(clknet_1_1__leaf__04680_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04682_ (.A(clknet_0__04682_),
    .X(clknet_1_1__leaf__04682_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04685_ (.A(clknet_0__04685_),
    .X(clknet_1_1__leaf__04685_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f__04686_ (.A(clknet_0__04686_),
    .X(clknet_1_1__leaf__04686_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_user_clock1 (.A(clknet_0_user_clock1),
    .X(clknet_1_1__leaf_user_clock1));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_user_clock2 (.A(clknet_0_user_clock2),
    .X(clknet_1_1__leaf_user_clock2));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_0_0_mclk (.A(net1695),
    .X(clknet_2_0_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04353_ (.A(clknet_0__04353_),
    .X(clknet_2_0__leaf__04353_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04358_ (.A(clknet_0__04358_),
    .X(clknet_2_0__leaf__04358_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04359_ (.A(clknet_0__04359_),
    .X(clknet_2_0__leaf__04359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04493_ (.A(clknet_0__04493_),
    .X(clknet_2_0__leaf__04493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04564_ (.A(clknet_0__04564_),
    .X(clknet_2_0__leaf__04564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04567_ (.A(clknet_0__04567_),
    .X(clknet_2_0__leaf__04567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04586_ (.A(clknet_0__04586_),
    .X(clknet_2_0__leaf__04586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04589_ (.A(clknet_0__04589_),
    .X(clknet_2_0__leaf__04589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04608_ (.A(clknet_0__04608_),
    .X(clknet_2_0__leaf__04608_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04611_ (.A(clknet_0__04611_),
    .X(clknet_2_0__leaf__04611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04633_ (.A(clknet_0__04633_),
    .X(clknet_2_0__leaf__04633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f__04653_ (.A(clknet_0__04653_),
    .X(clknet_2_0__leaf__04653_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_1_0_mclk (.A(clknet_0_mclk),
    .X(clknet_2_1_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04353_ (.A(clknet_0__04353_),
    .X(clknet_2_1__leaf__04353_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04358_ (.A(clknet_0__04358_),
    .X(clknet_2_1__leaf__04358_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04359_ (.A(clknet_0__04359_),
    .X(clknet_2_1__leaf__04359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04493_ (.A(clknet_0__04493_),
    .X(clknet_2_1__leaf__04493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04564_ (.A(clknet_0__04564_),
    .X(clknet_2_1__leaf__04564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04567_ (.A(clknet_0__04567_),
    .X(clknet_2_1__leaf__04567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04586_ (.A(clknet_0__04586_),
    .X(clknet_2_1__leaf__04586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04589_ (.A(clknet_0__04589_),
    .X(clknet_2_1__leaf__04589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04608_ (.A(clknet_0__04608_),
    .X(clknet_2_1__leaf__04608_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04611_ (.A(clknet_0__04611_),
    .X(clknet_2_1__leaf__04611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04633_ (.A(clknet_0__04633_),
    .X(clknet_2_1__leaf__04633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f__04653_ (.A(clknet_0__04653_),
    .X(clknet_2_1__leaf__04653_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_2_0_mclk (.A(net1696),
    .X(clknet_2_2_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04353_ (.A(clknet_0__04353_),
    .X(clknet_2_2__leaf__04353_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04358_ (.A(clknet_0__04358_),
    .X(clknet_2_2__leaf__04358_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04359_ (.A(clknet_0__04359_),
    .X(clknet_2_2__leaf__04359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04493_ (.A(clknet_0__04493_),
    .X(clknet_2_2__leaf__04493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04564_ (.A(clknet_0__04564_),
    .X(clknet_2_2__leaf__04564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04567_ (.A(clknet_0__04567_),
    .X(clknet_2_2__leaf__04567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04586_ (.A(clknet_0__04586_),
    .X(clknet_2_2__leaf__04586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04589_ (.A(clknet_0__04589_),
    .X(clknet_2_2__leaf__04589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04608_ (.A(clknet_0__04608_),
    .X(clknet_2_2__leaf__04608_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04611_ (.A(clknet_0__04611_),
    .X(clknet_2_2__leaf__04611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04633_ (.A(clknet_0__04633_),
    .X(clknet_2_2__leaf__04633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f__04653_ (.A(clknet_0__04653_),
    .X(clknet_2_2__leaf__04653_));
 sky130_fd_sc_hd__clkbuf_8 clkbuf_2_3_0_mclk (.A(net1696),
    .X(clknet_2_3_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04353_ (.A(clknet_0__04353_),
    .X(clknet_2_3__leaf__04353_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04358_ (.A(clknet_0__04358_),
    .X(clknet_2_3__leaf__04358_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04359_ (.A(clknet_0__04359_),
    .X(clknet_2_3__leaf__04359_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04493_ (.A(clknet_0__04493_),
    .X(clknet_2_3__leaf__04493_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04564_ (.A(clknet_0__04564_),
    .X(clknet_2_3__leaf__04564_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04567_ (.A(clknet_0__04567_),
    .X(clknet_2_3__leaf__04567_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04586_ (.A(clknet_0__04586_),
    .X(clknet_2_3__leaf__04586_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04589_ (.A(clknet_0__04589_),
    .X(clknet_2_3__leaf__04589_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04608_ (.A(clknet_0__04608_),
    .X(clknet_2_3__leaf__04608_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04611_ (.A(clknet_0__04611_),
    .X(clknet_2_3__leaf__04611_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04633_ (.A(clknet_0__04633_),
    .X(clknet_2_3__leaf__04633_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f__04653_ (.A(clknet_0__04653_),
    .X(clknet_2_3__leaf__04653_));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_0__f_mclk (.A(clknet_2_0_0_mclk),
    .X(clknet_4_0__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_10__f_mclk (.A(clknet_2_2_0_mclk),
    .X(clknet_4_10__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_11__f_mclk (.A(clknet_2_2_0_mclk),
    .X(clknet_4_11__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_12__f_mclk (.A(clknet_2_3_0_mclk),
    .X(clknet_4_12__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_13__f_mclk (.A(clknet_2_3_0_mclk),
    .X(clknet_4_13__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_14__f_mclk (.A(clknet_2_3_0_mclk),
    .X(clknet_4_14__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_15__f_mclk (.A(clknet_2_3_0_mclk),
    .X(clknet_4_15__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_1__f_mclk (.A(clknet_2_0_0_mclk),
    .X(clknet_4_1__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_2__f_mclk (.A(clknet_2_0_0_mclk),
    .X(clknet_4_2__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_3__f_mclk (.A(clknet_2_0_0_mclk),
    .X(clknet_4_3__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_4__f_mclk (.A(clknet_2_1_0_mclk),
    .X(clknet_4_4__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_5__f_mclk (.A(clknet_2_1_0_mclk),
    .X(clknet_4_5__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_6__f_mclk (.A(clknet_2_1_0_mclk),
    .X(clknet_4_6__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_7__f_mclk (.A(clknet_2_1_0_mclk),
    .X(clknet_4_7__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_8__f_mclk (.A(clknet_2_2_0_mclk),
    .X(clknet_4_8__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_4_9__f_mclk (.A(clknet_2_2_0_mclk),
    .X(clknet_4_9__leaf_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_0_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_0_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_100_mclk (.A(clknet_4_4__leaf_mclk),
    .X(clknet_leaf_100_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_102_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_102_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_103_mclk (.A(clknet_4_4__leaf_mclk),
    .X(clknet_leaf_103_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_104_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_104_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_105_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_105_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_106_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_106_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_107_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_107_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_109_mclk (.A(clknet_4_4__leaf_mclk),
    .X(clknet_leaf_109_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_10_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_10_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_110_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_110_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_111_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_111_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_112_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_112_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_113_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_113_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_114_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_114_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_115_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_115_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_116_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_116_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_117_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_117_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_118_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_118_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_11_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_11_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_120_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_120_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_122_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_122_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_123_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_123_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_124_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_124_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_126_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_126_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_127_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_127_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_128_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_128_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_12_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_12_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_13_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_13_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_14_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_14_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_15_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_15_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_16_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_16_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_17_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_17_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_19_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_19_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_1_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_1_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_20_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_20_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_21_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_21_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_22_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_22_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_23_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_23_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_24_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_24_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_25_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_25_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_26_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_26_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_28_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_28_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_29_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_29_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_2_mclk (.A(clknet_4_0__leaf_mclk),
    .X(clknet_leaf_2_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_30_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_30_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_31_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_31_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_32_mclk (.A(clknet_4_8__leaf_mclk),
    .X(clknet_leaf_32_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_33_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_33_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_34_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_34_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_35_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_35_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_36_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_36_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_37_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_37_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_38_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_38_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_39_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_39_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_40_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_40_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_41_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_41_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_42_mclk (.A(clknet_4_10__leaf_mclk),
    .X(clknet_leaf_42_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_43_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_43_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_44_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_44_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_45_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_45_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_46_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_46_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_47_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_47_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_48_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_48_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_4_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_4_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_51_mclk (.A(clknet_4_11__leaf_mclk),
    .X(clknet_leaf_51_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_53_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_53_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_54_mclk (.A(clknet_4_9__leaf_mclk),
    .X(clknet_leaf_54_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_55_mclk (.A(clknet_4_12__leaf_mclk),
    .X(clknet_leaf_55_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_56_mclk (.A(clknet_4_12__leaf_mclk),
    .X(clknet_leaf_56_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_58_mclk (.A(clknet_4_12__leaf_mclk),
    .X(clknet_leaf_58_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_5_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_5_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_60_mclk (.A(clknet_4_14__leaf_mclk),
    .X(clknet_leaf_60_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_62_mclk (.A(clknet_4_15__leaf_mclk),
    .X(clknet_leaf_62_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_63_mclk (.A(clknet_4_14__leaf_mclk),
    .X(clknet_leaf_63_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_65_mclk (.A(clknet_4_14__leaf_mclk),
    .X(clknet_leaf_65_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_66_mclk (.A(clknet_4_15__leaf_mclk),
    .X(clknet_leaf_66_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_67_mclk (.A(clknet_4_15__leaf_mclk),
    .X(clknet_leaf_67_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_69_mclk (.A(clknet_4_15__leaf_mclk),
    .X(clknet_leaf_69_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_6_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_6_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_70_mclk (.A(clknet_4_15__leaf_mclk),
    .X(clknet_leaf_70_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_72_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_72_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_73_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_73_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_74_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_74_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_75_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_75_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_76_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_76_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_77_mclk (.A(clknet_4_13__leaf_mclk),
    .X(clknet_leaf_77_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_78_mclk (.A(clknet_4_12__leaf_mclk),
    .X(clknet_leaf_78_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_79_mclk (.A(clknet_4_12__leaf_mclk),
    .X(clknet_leaf_79_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_7_mclk (.A(clknet_4_2__leaf_mclk),
    .X(clknet_leaf_7_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_80_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_80_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_81_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_81_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_82_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_82_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_83_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_83_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_84_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_84_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_85_mclk (.A(clknet_4_6__leaf_mclk),
    .X(clknet_leaf_85_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_86_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_86_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_87_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_87_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_88_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_88_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_89_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_89_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_8_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_8_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_90_mclk (.A(clknet_4_7__leaf_mclk),
    .X(clknet_leaf_90_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_91_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_91_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_92_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_92_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_93_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_93_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_94_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_94_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_95_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_95_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_96_mclk (.A(clknet_4_5__leaf_mclk),
    .X(clknet_leaf_96_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_97_mclk (.A(clknet_4_4__leaf_mclk),
    .X(clknet_leaf_97_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_99_mclk (.A(clknet_4_1__leaf_mclk),
    .X(clknet_leaf_99_mclk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_leaf_9_mclk (.A(clknet_4_3__leaf_mclk),
    .X(clknet_leaf_9_mclk));
 sky130_fd_sc_hd__clkbuf_4 fanout1000 (.A(net1002),
    .X(net1000));
 sky130_fd_sc_hd__clkbuf_2 fanout1001 (.A(net1002),
    .X(net1001));
 sky130_fd_sc_hd__clkbuf_2 fanout1002 (.A(net1011),
    .X(net1002));
 sky130_fd_sc_hd__clkbuf_4 fanout1003 (.A(net1006),
    .X(net1003));
 sky130_fd_sc_hd__clkbuf_4 fanout1004 (.A(net1006),
    .X(net1004));
 sky130_fd_sc_hd__buf_2 fanout1005 (.A(net1006),
    .X(net1005));
 sky130_fd_sc_hd__clkbuf_2 fanout1006 (.A(net1011),
    .X(net1006));
 sky130_fd_sc_hd__clkbuf_4 fanout1007 (.A(net1011),
    .X(net1007));
 sky130_fd_sc_hd__clkbuf_4 fanout1008 (.A(net1010),
    .X(net1008));
 sky130_fd_sc_hd__clkbuf_2 fanout1009 (.A(net1010),
    .X(net1009));
 sky130_fd_sc_hd__buf_2 fanout1010 (.A(net1011),
    .X(net1010));
 sky130_fd_sc_hd__buf_2 fanout1011 (.A(net1041),
    .X(net1011));
 sky130_fd_sc_hd__clkbuf_4 fanout1012 (.A(net1013),
    .X(net1012));
 sky130_fd_sc_hd__clkbuf_2 fanout1013 (.A(net1017),
    .X(net1013));
 sky130_fd_sc_hd__clkbuf_4 fanout1014 (.A(net1015),
    .X(net1014));
 sky130_fd_sc_hd__clkbuf_4 fanout1015 (.A(net1016),
    .X(net1015));
 sky130_fd_sc_hd__buf_2 fanout1016 (.A(net1017),
    .X(net1016));
 sky130_fd_sc_hd__clkbuf_2 fanout1017 (.A(net1041),
    .X(net1017));
 sky130_fd_sc_hd__clkbuf_4 fanout1018 (.A(net1023),
    .X(net1018));
 sky130_fd_sc_hd__clkbuf_4 fanout1019 (.A(net1020),
    .X(net1019));
 sky130_fd_sc_hd__buf_2 fanout1020 (.A(net1023),
    .X(net1020));
 sky130_fd_sc_hd__buf_4 fanout1021 (.A(net1022),
    .X(net1021));
 sky130_fd_sc_hd__buf_4 fanout1022 (.A(net1023),
    .X(net1022));
 sky130_fd_sc_hd__clkbuf_4 fanout1023 (.A(net1041),
    .X(net1023));
 sky130_fd_sc_hd__clkbuf_4 fanout1024 (.A(net1025),
    .X(net1024));
 sky130_fd_sc_hd__clkbuf_4 fanout1025 (.A(net1030),
    .X(net1025));
 sky130_fd_sc_hd__clkbuf_4 fanout1026 (.A(net1027),
    .X(net1026));
 sky130_fd_sc_hd__clkbuf_4 fanout1027 (.A(net1030),
    .X(net1027));
 sky130_fd_sc_hd__clkbuf_4 fanout1028 (.A(net1030),
    .X(net1028));
 sky130_fd_sc_hd__clkbuf_4 fanout1029 (.A(net1030),
    .X(net1029));
 sky130_fd_sc_hd__buf_2 fanout1030 (.A(net1041),
    .X(net1030));
 sky130_fd_sc_hd__clkbuf_4 fanout1031 (.A(net1035),
    .X(net1031));
 sky130_fd_sc_hd__buf_2 fanout1032 (.A(net1035),
    .X(net1032));
 sky130_fd_sc_hd__clkbuf_4 fanout1033 (.A(net1034),
    .X(net1033));
 sky130_fd_sc_hd__clkbuf_4 fanout1034 (.A(net1035),
    .X(net1034));
 sky130_fd_sc_hd__clkbuf_4 fanout1035 (.A(net1040),
    .X(net1035));
 sky130_fd_sc_hd__buf_4 fanout1036 (.A(net1038),
    .X(net1036));
 sky130_fd_sc_hd__buf_2 fanout1037 (.A(net1038),
    .X(net1037));
 sky130_fd_sc_hd__clkbuf_4 fanout1038 (.A(net1039),
    .X(net1038));
 sky130_fd_sc_hd__clkbuf_4 fanout1039 (.A(net1040),
    .X(net1039));
 sky130_fd_sc_hd__buf_2 fanout1040 (.A(net1041),
    .X(net1040));
 sky130_fd_sc_hd__buf_6 fanout1041 (.A(net1043),
    .X(net1041));
 sky130_fd_sc_hd__buf_6 fanout1042 (.A(\u_glbl_reg.s_reset_n ),
    .X(net1042));
 sky130_fd_sc_hd__clkbuf_4 fanout1044 (.A(net1045),
    .X(net1044));
 sky130_fd_sc_hd__clkbuf_4 fanout1045 (.A(net1061),
    .X(net1045));
 sky130_fd_sc_hd__clkbuf_4 fanout1046 (.A(net1047),
    .X(net1046));
 sky130_fd_sc_hd__buf_2 fanout1047 (.A(net1061),
    .X(net1047));
 sky130_fd_sc_hd__clkbuf_4 fanout1048 (.A(net1049),
    .X(net1048));
 sky130_fd_sc_hd__clkbuf_4 fanout1049 (.A(net1051),
    .X(net1049));
 sky130_fd_sc_hd__clkbuf_4 fanout1050 (.A(net1051),
    .X(net1050));
 sky130_fd_sc_hd__clkbuf_2 fanout1051 (.A(net1061),
    .X(net1051));
 sky130_fd_sc_hd__clkbuf_4 fanout1052 (.A(net1054),
    .X(net1052));
 sky130_fd_sc_hd__clkbuf_2 fanout1053 (.A(net1054),
    .X(net1053));
 sky130_fd_sc_hd__clkbuf_4 fanout1054 (.A(net1061),
    .X(net1054));
 sky130_fd_sc_hd__clkbuf_4 fanout1055 (.A(net1057),
    .X(net1055));
 sky130_fd_sc_hd__clkbuf_4 fanout1056 (.A(net1057),
    .X(net1056));
 sky130_fd_sc_hd__clkbuf_4 fanout1057 (.A(net1061),
    .X(net1057));
 sky130_fd_sc_hd__buf_4 fanout1058 (.A(net1060),
    .X(net1058));
 sky130_fd_sc_hd__buf_4 fanout1059 (.A(net1060),
    .X(net1059));
 sky130_fd_sc_hd__clkbuf_4 fanout1060 (.A(net1061),
    .X(net1060));
 sky130_fd_sc_hd__buf_4 fanout1061 (.A(net1068),
    .X(net1061));
 sky130_fd_sc_hd__buf_4 fanout1062 (.A(net1063),
    .X(net1062));
 sky130_fd_sc_hd__buf_4 fanout1063 (.A(net1069),
    .X(net1063));
 sky130_fd_sc_hd__clkbuf_4 fanout1064 (.A(net1066),
    .X(net1064));
 sky130_fd_sc_hd__clkbuf_2 fanout1065 (.A(net1066),
    .X(net1065));
 sky130_fd_sc_hd__clkbuf_4 fanout1066 (.A(net1067),
    .X(net1066));
 sky130_fd_sc_hd__clkbuf_4 fanout1067 (.A(net1069),
    .X(net1067));
 sky130_fd_sc_hd__buf_6 fanout1068 (.A(\u_glbl_reg.p_reset_n ),
    .X(net1068));
 sky130_fd_sc_hd__buf_12 fanout1070 (.A(net1071),
    .X(net1070));
 sky130_fd_sc_hd__buf_12 fanout1071 (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[15] ),
    .X(net1071));
 sky130_fd_sc_hd__buf_4 fanout1072 (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[14] ),
    .X(net1072));
 sky130_fd_sc_hd__buf_4 fanout1073 (.A(\u_pwm.u_pwm_2.u_pwm.pwm_cnt[10] ),
    .X(net1073));
 sky130_fd_sc_hd__buf_12 fanout1074 (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ),
    .X(net1074));
 sky130_fd_sc_hd__buf_8 fanout1075 (.A(\u_pwm.u_pwm_1.u_pwm.pwm_cnt[15] ),
    .X(net1075));
 sky130_fd_sc_hd__buf_12 fanout1076 (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[15] ),
    .X(net1076));
 sky130_fd_sc_hd__buf_8 fanout1077 (.A(\u_pwm.u_pwm_0.u_pwm.pwm_cnt[15] ),
    .X(net1077));
 sky130_fd_sc_hd__buf_4 fanout1080 (.A(net1082),
    .X(net1080));
 sky130_fd_sc_hd__clkbuf_4 fanout1081 (.A(net1082),
    .X(net1081));
 sky130_fd_sc_hd__clkbuf_4 fanout1082 (.A(\u_ws281x.u_reg.gfifo[0].u_fifo.rd_ptr ),
    .X(net1082));
 sky130_fd_sc_hd__buf_4 fanout1083 (.A(net1085),
    .X(net1083));
 sky130_fd_sc_hd__buf_4 fanout1084 (.A(net1085),
    .X(net1084));
 sky130_fd_sc_hd__clkbuf_4 fanout1085 (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.rd_ptr ),
    .X(net1085));
 sky130_fd_sc_hd__buf_2 fanout1086 (.A(net1090),
    .X(net1086));
 sky130_fd_sc_hd__clkbuf_2 fanout1087 (.A(net1090),
    .X(net1087));
 sky130_fd_sc_hd__clkbuf_4 fanout1088 (.A(net1090),
    .X(net1088));
 sky130_fd_sc_hd__clkbuf_2 fanout1089 (.A(net1090),
    .X(net1089));
 sky130_fd_sc_hd__clkbuf_4 fanout1090 (.A(\reg_blk_sel[3] ),
    .X(net1090));
 sky130_fd_sc_hd__clkbuf_4 fanout1091 (.A(\reg_blk_sel[0] ),
    .X(net1091));
 sky130_fd_sc_hd__buf_2 fanout1092 (.A(\reg_blk_sel[0] ),
    .X(net1092));
 sky130_fd_sc_hd__buf_6 fanout1109 (.A(\u_glbl_reg.cfg_multi_func_sel[30] ),
    .X(net1109));
 sky130_fd_sc_hd__clkbuf_4 fanout1110 (.A(_03462_),
    .X(net1110));
 sky130_fd_sc_hd__buf_2 fanout1111 (.A(net1112),
    .X(net1111));
 sky130_fd_sc_hd__buf_2 fanout1112 (.A(net1113),
    .X(net1112));
 sky130_fd_sc_hd__buf_2 fanout1113 (.A(_03460_),
    .X(net1113));
 sky130_fd_sc_hd__buf_2 fanout1114 (.A(net1115),
    .X(net1114));
 sky130_fd_sc_hd__buf_2 fanout1115 (.A(net1118),
    .X(net1115));
 sky130_fd_sc_hd__clkbuf_4 fanout1116 (.A(net1117),
    .X(net1116));
 sky130_fd_sc_hd__buf_2 fanout1117 (.A(net1118),
    .X(net1117));
 sky130_fd_sc_hd__buf_2 fanout1118 (.A(_03457_),
    .X(net1118));
 sky130_fd_sc_hd__buf_2 fanout1119 (.A(net1120),
    .X(net1119));
 sky130_fd_sc_hd__buf_2 fanout1120 (.A(net1123),
    .X(net1120));
 sky130_fd_sc_hd__clkbuf_4 fanout1121 (.A(net1122),
    .X(net1121));
 sky130_fd_sc_hd__buf_2 fanout1122 (.A(net1123),
    .X(net1122));
 sky130_fd_sc_hd__buf_2 fanout1123 (.A(_03456_),
    .X(net1123));
 sky130_fd_sc_hd__buf_4 fanout1124 (.A(net1126),
    .X(net1124));
 sky130_fd_sc_hd__clkbuf_2 fanout1125 (.A(net1126),
    .X(net1125));
 sky130_fd_sc_hd__buf_2 fanout1126 (.A(_01546_),
    .X(net1126));
 sky130_fd_sc_hd__clkbuf_4 fanout1127 (.A(net1128),
    .X(net1127));
 sky130_fd_sc_hd__clkbuf_2 fanout1128 (.A(_01546_),
    .X(net1128));
 sky130_fd_sc_hd__buf_2 fanout1129 (.A(_01543_),
    .X(net1129));
 sky130_fd_sc_hd__clkbuf_2 fanout1130 (.A(_01543_),
    .X(net1130));
 sky130_fd_sc_hd__clkbuf_4 fanout1131 (.A(net1132),
    .X(net1131));
 sky130_fd_sc_hd__buf_4 fanout1132 (.A(net1133),
    .X(net1132));
 sky130_fd_sc_hd__buf_4 fanout1133 (.A(_01541_),
    .X(net1133));
 sky130_fd_sc_hd__buf_4 fanout1134 (.A(_01541_),
    .X(net1134));
 sky130_fd_sc_hd__clkbuf_4 fanout1135 (.A(_01541_),
    .X(net1135));
 sky130_fd_sc_hd__clkbuf_4 fanout1136 (.A(net1141),
    .X(net1136));
 sky130_fd_sc_hd__buf_2 fanout1137 (.A(net1141),
    .X(net1137));
 sky130_fd_sc_hd__buf_4 fanout1138 (.A(net1141),
    .X(net1138));
 sky130_fd_sc_hd__clkbuf_4 fanout1139 (.A(net1140),
    .X(net1139));
 sky130_fd_sc_hd__buf_4 fanout1140 (.A(net1141),
    .X(net1140));
 sky130_fd_sc_hd__clkbuf_4 fanout1141 (.A(_01540_),
    .X(net1141));
 sky130_fd_sc_hd__buf_4 fanout1142 (.A(net1144),
    .X(net1142));
 sky130_fd_sc_hd__buf_4 fanout1143 (.A(net1144),
    .X(net1143));
 sky130_fd_sc_hd__buf_4 fanout1144 (.A(_01349_),
    .X(net1144));
 sky130_fd_sc_hd__buf_4 fanout1145 (.A(net1147),
    .X(net1145));
 sky130_fd_sc_hd__clkbuf_2 fanout1146 (.A(net1147),
    .X(net1146));
 sky130_fd_sc_hd__clkbuf_8 fanout1147 (.A(net1151),
    .X(net1147));
 sky130_fd_sc_hd__buf_2 fanout1148 (.A(net1149),
    .X(net1148));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1149 (.A(net1151),
    .X(net1149));
 sky130_fd_sc_hd__clkbuf_4 fanout1150 (.A(net1151),
    .X(net1150));
 sky130_fd_sc_hd__buf_4 fanout1151 (.A(_01349_),
    .X(net1151));
 sky130_fd_sc_hd__buf_2 fanout1152 (.A(net1153),
    .X(net1152));
 sky130_fd_sc_hd__buf_2 fanout1153 (.A(_01116_),
    .X(net1153));
 sky130_fd_sc_hd__clkbuf_4 fanout1154 (.A(net1159),
    .X(net1154));
 sky130_fd_sc_hd__clkbuf_4 fanout1155 (.A(net1159),
    .X(net1155));
 sky130_fd_sc_hd__buf_2 fanout1156 (.A(net1159),
    .X(net1156));
 sky130_fd_sc_hd__buf_4 fanout1157 (.A(net1159),
    .X(net1157));
 sky130_fd_sc_hd__clkbuf_4 fanout1158 (.A(net1159),
    .X(net1158));
 sky130_fd_sc_hd__buf_4 fanout1159 (.A(_01114_),
    .X(net1159));
 sky130_fd_sc_hd__clkbuf_4 fanout1160 (.A(net1161),
    .X(net1160));
 sky130_fd_sc_hd__clkbuf_4 fanout1161 (.A(_01114_),
    .X(net1161));
 sky130_fd_sc_hd__clkbuf_4 fanout1162 (.A(net1163),
    .X(net1162));
 sky130_fd_sc_hd__buf_4 fanout1163 (.A(_01114_),
    .X(net1163));
 sky130_fd_sc_hd__clkbuf_2 fanout1164 (.A(net1165),
    .X(net1164));
 sky130_fd_sc_hd__clkbuf_4 fanout1165 (.A(_01114_),
    .X(net1165));
 sky130_fd_sc_hd__buf_2 fanout1166 (.A(net1171),
    .X(net1166));
 sky130_fd_sc_hd__buf_2 fanout1167 (.A(net1171),
    .X(net1167));
 sky130_fd_sc_hd__buf_2 fanout1168 (.A(net1171),
    .X(net1168));
 sky130_fd_sc_hd__buf_2 fanout1169 (.A(net1170),
    .X(net1169));
 sky130_fd_sc_hd__buf_4 fanout1170 (.A(net1171),
    .X(net1170));
 sky130_fd_sc_hd__clkbuf_4 fanout1171 (.A(_01113_),
    .X(net1171));
 sky130_fd_sc_hd__clkbuf_4 fanout1172 (.A(net1174),
    .X(net1172));
 sky130_fd_sc_hd__clkbuf_2 fanout1173 (.A(net1174),
    .X(net1173));
 sky130_fd_sc_hd__buf_4 fanout1174 (.A(_01113_),
    .X(net1174));
 sky130_fd_sc_hd__buf_2 fanout1175 (.A(net1178),
    .X(net1175));
 sky130_fd_sc_hd__clkbuf_2 fanout1176 (.A(net1178),
    .X(net1176));
 sky130_fd_sc_hd__buf_4 fanout1177 (.A(net1178),
    .X(net1177));
 sky130_fd_sc_hd__buf_2 fanout1178 (.A(_01004_),
    .X(net1178));
 sky130_fd_sc_hd__buf_4 fanout1179 (.A(_00998_),
    .X(net1179));
 sky130_fd_sc_hd__clkbuf_4 fanout1180 (.A(_00998_),
    .X(net1180));
 sky130_fd_sc_hd__clkbuf_4 fanout1181 (.A(net1182),
    .X(net1181));
 sky130_fd_sc_hd__clkbuf_4 fanout1182 (.A(_00996_),
    .X(net1182));
 sky130_fd_sc_hd__clkbuf_2 fanout1201 (.A(net1202),
    .X(net1201));
 sky130_fd_sc_hd__buf_2 fanout1202 (.A(net2293),
    .X(net1202));
 sky130_fd_sc_hd__buf_2 fanout1203 (.A(net1205),
    .X(net1203));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1204 (.A(net1205),
    .X(net1204));
 sky130_fd_sc_hd__clkbuf_2 fanout1205 (.A(net2293),
    .X(net1205));
 sky130_fd_sc_hd__clkbuf_4 fanout1207 (.A(net1208),
    .X(net1207));
 sky130_fd_sc_hd__clkbuf_2 fanout1208 (.A(net1209),
    .X(net1208));
 sky130_fd_sc_hd__buf_4 fanout1209 (.A(net1729),
    .X(net1209));
 sky130_fd_sc_hd__buf_4 fanout1210 (.A(net1729),
    .X(net1210));
 sky130_fd_sc_hd__clkbuf_8 fanout1211 (.A(net1213),
    .X(net1211));
 sky130_fd_sc_hd__buf_6 fanout1212 (.A(net1213),
    .X(net1212));
 sky130_fd_sc_hd__clkbuf_8 fanout1213 (.A(_01350_),
    .X(net1213));
 sky130_fd_sc_hd__clkbuf_4 fanout1214 (.A(net1216),
    .X(net1214));
 sky130_fd_sc_hd__buf_2 fanout1215 (.A(net1216),
    .X(net1215));
 sky130_fd_sc_hd__clkbuf_4 fanout1216 (.A(_01129_),
    .X(net1216));
 sky130_fd_sc_hd__clkbuf_4 fanout1217 (.A(net1218),
    .X(net1217));
 sky130_fd_sc_hd__clkbuf_4 fanout1218 (.A(net1221),
    .X(net1218));
 sky130_fd_sc_hd__clkbuf_4 fanout1219 (.A(net1220),
    .X(net1219));
 sky130_fd_sc_hd__buf_4 fanout1220 (.A(net1221),
    .X(net1220));
 sky130_fd_sc_hd__clkbuf_4 fanout1221 (.A(net1225),
    .X(net1221));
 sky130_fd_sc_hd__buf_4 fanout1222 (.A(net1225),
    .X(net1222));
 sky130_fd_sc_hd__clkbuf_4 fanout1223 (.A(net1224),
    .X(net1223));
 sky130_fd_sc_hd__clkbuf_4 fanout1224 (.A(net1225),
    .X(net1224));
 sky130_fd_sc_hd__clkbuf_4 fanout1225 (.A(_01007_),
    .X(net1225));
 sky130_fd_sc_hd__clkbuf_4 fanout1226 (.A(net1227),
    .X(net1226));
 sky130_fd_sc_hd__buf_2 fanout1227 (.A(net1228),
    .X(net1227));
 sky130_fd_sc_hd__clkbuf_4 fanout1228 (.A(net1233),
    .X(net1228));
 sky130_fd_sc_hd__clkbuf_4 fanout1229 (.A(net1230),
    .X(net1229));
 sky130_fd_sc_hd__buf_4 fanout1230 (.A(net1233),
    .X(net1230));
 sky130_fd_sc_hd__buf_2 fanout1231 (.A(net1233),
    .X(net1231));
 sky130_fd_sc_hd__clkbuf_4 fanout1232 (.A(net1233),
    .X(net1232));
 sky130_fd_sc_hd__buf_4 fanout1233 (.A(_01007_),
    .X(net1233));
 sky130_fd_sc_hd__clkbuf_4 fanout1234 (.A(net1235),
    .X(net1234));
 sky130_fd_sc_hd__buf_2 fanout1235 (.A(net1253),
    .X(net1235));
 sky130_fd_sc_hd__clkbuf_4 fanout1236 (.A(net1238),
    .X(net1236));
 sky130_fd_sc_hd__clkbuf_4 fanout1237 (.A(net1238),
    .X(net1237));
 sky130_fd_sc_hd__clkbuf_4 fanout1238 (.A(net1253),
    .X(net1238));
 sky130_fd_sc_hd__clkbuf_4 fanout1239 (.A(net1242),
    .X(net1239));
 sky130_fd_sc_hd__clkbuf_2 fanout1240 (.A(net1242),
    .X(net1240));
 sky130_fd_sc_hd__clkbuf_4 fanout1241 (.A(net1242),
    .X(net1241));
 sky130_fd_sc_hd__clkbuf_4 fanout1242 (.A(net1253),
    .X(net1242));
 sky130_fd_sc_hd__clkbuf_4 fanout1243 (.A(net1247),
    .X(net1243));
 sky130_fd_sc_hd__clkbuf_2 fanout1244 (.A(net1247),
    .X(net1244));
 sky130_fd_sc_hd__clkbuf_4 fanout1245 (.A(net1247),
    .X(net1245));
 sky130_fd_sc_hd__clkbuf_2 fanout1246 (.A(net1247),
    .X(net1246));
 sky130_fd_sc_hd__buf_4 fanout1247 (.A(net1253),
    .X(net1247));
 sky130_fd_sc_hd__clkbuf_4 fanout1248 (.A(net1252),
    .X(net1248));
 sky130_fd_sc_hd__clkbuf_2 fanout1249 (.A(net1252),
    .X(net1249));
 sky130_fd_sc_hd__buf_2 fanout1250 (.A(net1251),
    .X(net1250));
 sky130_fd_sc_hd__clkbuf_2 fanout1251 (.A(net1252),
    .X(net1251));
 sky130_fd_sc_hd__clkbuf_2 fanout1252 (.A(net1253),
    .X(net1252));
 sky130_fd_sc_hd__clkbuf_4 fanout1253 (.A(_01006_),
    .X(net1253));
 sky130_fd_sc_hd__clkbuf_2 fanout1254 (.A(net1255),
    .X(net1254));
 sky130_fd_sc_hd__clkbuf_4 fanout1255 (.A(_00794_),
    .X(net1255));
 sky130_fd_sc_hd__clkbuf_4 fanout1256 (.A(net1257),
    .X(net1256));
 sky130_fd_sc_hd__clkbuf_4 fanout1257 (.A(net1259),
    .X(net1257));
 sky130_fd_sc_hd__buf_4 fanout1258 (.A(net1259),
    .X(net1258));
 sky130_fd_sc_hd__clkbuf_4 fanout1259 (.A(net1265),
    .X(net1259));
 sky130_fd_sc_hd__buf_6 fanout1260 (.A(net1265),
    .X(net1260));
 sky130_fd_sc_hd__clkbuf_4 fanout1261 (.A(net1265),
    .X(net1261));
 sky130_fd_sc_hd__clkbuf_4 fanout1262 (.A(net1264),
    .X(net1262));
 sky130_fd_sc_hd__buf_2 fanout1263 (.A(net1264),
    .X(net1263));
 sky130_fd_sc_hd__clkbuf_4 fanout1264 (.A(net1265),
    .X(net1264));
 sky130_fd_sc_hd__clkbuf_4 fanout1265 (.A(_00778_),
    .X(net1265));
 sky130_fd_sc_hd__clkbuf_4 fanout1266 (.A(net1267),
    .X(net1266));
 sky130_fd_sc_hd__clkbuf_8 fanout1267 (.A(net1270),
    .X(net1267));
 sky130_fd_sc_hd__clkbuf_4 fanout1268 (.A(net1269),
    .X(net1268));
 sky130_fd_sc_hd__buf_4 fanout1269 (.A(net1270),
    .X(net1269));
 sky130_fd_sc_hd__clkbuf_4 fanout1270 (.A(net1284),
    .X(net1270));
 sky130_fd_sc_hd__buf_6 fanout1271 (.A(net1284),
    .X(net1271));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1272 (.A(net1285),
    .X(net1272));
 sky130_fd_sc_hd__clkbuf_4 fanout1273 (.A(net1274),
    .X(net1273));
 sky130_fd_sc_hd__clkbuf_4 fanout1274 (.A(net1284),
    .X(net1274));
 sky130_fd_sc_hd__buf_2 fanout1275 (.A(net1277),
    .X(net1275));
 sky130_fd_sc_hd__clkbuf_2 fanout1276 (.A(net1277),
    .X(net1276));
 sky130_fd_sc_hd__clkbuf_4 fanout1277 (.A(net1285),
    .X(net1277));
 sky130_fd_sc_hd__clkbuf_4 fanout1278 (.A(net1279),
    .X(net1278));
 sky130_fd_sc_hd__clkbuf_4 fanout1279 (.A(net1285),
    .X(net1279));
 sky130_fd_sc_hd__buf_2 fanout1280 (.A(net1283),
    .X(net1280));
 sky130_fd_sc_hd__clkbuf_2 fanout1281 (.A(net1283),
    .X(net1281));
 sky130_fd_sc_hd__clkbuf_2 fanout1282 (.A(net1283),
    .X(net1282));
 sky130_fd_sc_hd__buf_2 fanout1283 (.A(net1285),
    .X(net1283));
 sky130_fd_sc_hd__buf_6 fanout1284 (.A(_00777_),
    .X(net1284));
 sky130_fd_sc_hd__clkbuf_4 fanout1286 (.A(net1288),
    .X(net1286));
 sky130_fd_sc_hd__buf_2 fanout1287 (.A(net1288),
    .X(net1287));
 sky130_fd_sc_hd__clkbuf_4 fanout1288 (.A(net1290),
    .X(net1288));
 sky130_fd_sc_hd__clkbuf_8 fanout1289 (.A(net1290),
    .X(net1289));
 sky130_fd_sc_hd__buf_4 fanout1290 (.A(net99),
    .X(net1290));
 sky130_fd_sc_hd__buf_4 fanout1291 (.A(net1292),
    .X(net1291));
 sky130_fd_sc_hd__clkbuf_4 fanout1293 (.A(net1295),
    .X(net1293));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1294 (.A(net1295),
    .X(net1294));
 sky130_fd_sc_hd__clkbuf_4 fanout1295 (.A(net1298),
    .X(net1295));
 sky130_fd_sc_hd__clkbuf_4 fanout1296 (.A(net1298),
    .X(net1296));
 sky130_fd_sc_hd__clkbuf_2 fanout1297 (.A(net1298),
    .X(net1297));
 sky130_fd_sc_hd__buf_4 fanout1298 (.A(net98),
    .X(net1298));
 sky130_fd_sc_hd__buf_2 fanout1299 (.A(net1301),
    .X(net1299));
 sky130_fd_sc_hd__clkbuf_4 fanout1300 (.A(net1301),
    .X(net1300));
 sky130_fd_sc_hd__clkbuf_4 fanout1301 (.A(net1303),
    .X(net1301));
 sky130_fd_sc_hd__clkbuf_8 fanout1302 (.A(net1303),
    .X(net1302));
 sky130_fd_sc_hd__buf_4 fanout1303 (.A(net98),
    .X(net1303));
 sky130_fd_sc_hd__buf_2 fanout1308 (.A(net1311),
    .X(net1308));
 sky130_fd_sc_hd__clkbuf_2 fanout1309 (.A(net1311),
    .X(net1309));
 sky130_fd_sc_hd__clkbuf_4 fanout1310 (.A(net1311),
    .X(net1310));
 sky130_fd_sc_hd__buf_6 fanout1311 (.A(net1312),
    .X(net1311));
 sky130_fd_sc_hd__buf_6 fanout1312 (.A(net63),
    .X(net1312));
 sky130_fd_sc_hd__buf_4 fanout1316 (.A(net1317),
    .X(net1316));
 sky130_fd_sc_hd__buf_6 fanout1317 (.A(net62),
    .X(net1317));
 sky130_fd_sc_hd__clkbuf_4 fanout1319 (.A(net1320),
    .X(net1319));
 sky130_fd_sc_hd__clkbuf_4 fanout1320 (.A(net1321),
    .X(net1320));
 sky130_fd_sc_hd__buf_6 fanout1321 (.A(net62),
    .X(net1321));
 sky130_fd_sc_hd__clkbuf_4 fanout1323 (.A(net1325),
    .X(net1323));
 sky130_fd_sc_hd__buf_4 fanout1324 (.A(net1328),
    .X(net1324));
 sky130_fd_sc_hd__clkbuf_2 fanout1325 (.A(net1328),
    .X(net1325));
 sky130_fd_sc_hd__buf_6 fanout1326 (.A(net1328),
    .X(net1326));
 sky130_fd_sc_hd__buf_4 fanout1328 (.A(net61),
    .X(net1328));
 sky130_fd_sc_hd__buf_6 fanout1329 (.A(net1330),
    .X(net1329));
 sky130_fd_sc_hd__buf_2 fanout1331 (.A(net1332),
    .X(net1331));
 sky130_fd_sc_hd__clkbuf_4 fanout1332 (.A(net1333),
    .X(net1332));
 sky130_fd_sc_hd__clkbuf_4 fanout1333 (.A(net1338),
    .X(net1333));
 sky130_fd_sc_hd__clkbuf_4 fanout1334 (.A(net1335),
    .X(net1334));
 sky130_fd_sc_hd__buf_4 fanout1335 (.A(net1338),
    .X(net1335));
 sky130_fd_sc_hd__buf_6 fanout1336 (.A(net1338),
    .X(net1336));
 sky130_fd_sc_hd__buf_4 fanout1337 (.A(net1338),
    .X(net1337));
 sky130_fd_sc_hd__buf_4 fanout1343 (.A(net56),
    .X(net1343));
 sky130_fd_sc_hd__buf_2 fanout1344 (.A(net56),
    .X(net1344));
 sky130_fd_sc_hd__buf_4 fanout1346 (.A(net1347),
    .X(net1346));
 sky130_fd_sc_hd__buf_2 fanout1348 (.A(net1353),
    .X(net1348));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1349 (.A(net1353),
    .X(net1349));
 sky130_fd_sc_hd__buf_2 fanout1350 (.A(net1351),
    .X(net1350));
 sky130_fd_sc_hd__clkbuf_2 fanout1351 (.A(net1353),
    .X(net1351));
 sky130_fd_sc_hd__buf_2 fanout1352 (.A(net1353),
    .X(net1352));
 sky130_fd_sc_hd__buf_2 fanout1353 (.A(net53),
    .X(net1353));
 sky130_fd_sc_hd__buf_2 fanout1354 (.A(net1356),
    .X(net1354));
 sky130_fd_sc_hd__buf_2 fanout1355 (.A(net1356),
    .X(net1355));
 sky130_fd_sc_hd__buf_4 fanout1356 (.A(net1361),
    .X(net1356));
 sky130_fd_sc_hd__clkbuf_4 fanout1357 (.A(net1359),
    .X(net1357));
 sky130_fd_sc_hd__clkbuf_2 fanout1358 (.A(net1359),
    .X(net1358));
 sky130_fd_sc_hd__clkbuf_4 fanout1359 (.A(net1361),
    .X(net1359));
 sky130_fd_sc_hd__clkbuf_4 fanout1360 (.A(net1361),
    .X(net1360));
 sky130_fd_sc_hd__clkbuf_4 fanout1361 (.A(net53),
    .X(net1361));
 sky130_fd_sc_hd__buf_4 fanout1362 (.A(net1363),
    .X(net1362));
 sky130_fd_sc_hd__buf_4 fanout1363 (.A(net1364),
    .X(net1363));
 sky130_fd_sc_hd__buf_6 fanout1364 (.A(net1372),
    .X(net1364));
 sky130_fd_sc_hd__clkbuf_4 fanout1365 (.A(net1366),
    .X(net1365));
 sky130_fd_sc_hd__clkbuf_4 fanout1366 (.A(net1368),
    .X(net1366));
 sky130_fd_sc_hd__clkbuf_4 fanout1367 (.A(net1368),
    .X(net1367));
 sky130_fd_sc_hd__clkbuf_4 fanout1368 (.A(net1372),
    .X(net1368));
 sky130_fd_sc_hd__buf_2 fanout1369 (.A(net1371),
    .X(net1369));
 sky130_fd_sc_hd__clkbuf_2 fanout1370 (.A(net1371),
    .X(net1370));
 sky130_fd_sc_hd__clkbuf_2 fanout1371 (.A(net1372),
    .X(net1371));
 sky130_fd_sc_hd__buf_6 fanout1372 (.A(net52),
    .X(net1372));
 sky130_fd_sc_hd__clkbuf_4 fanout1378 (.A(net1383),
    .X(net1378));
 sky130_fd_sc_hd__buf_2 fanout1379 (.A(net1383),
    .X(net1379));
 sky130_fd_sc_hd__clkbuf_4 fanout1380 (.A(net1381),
    .X(net1380));
 sky130_fd_sc_hd__clkbuf_4 fanout1381 (.A(net1383),
    .X(net1381));
 sky130_fd_sc_hd__buf_4 fanout1382 (.A(net1383),
    .X(net1382));
 sky130_fd_sc_hd__clkbuf_4 fanout1383 (.A(net1384),
    .X(net1383));
 sky130_fd_sc_hd__clkbuf_4 fanout1384 (.A(net1385),
    .X(net1384));
 sky130_fd_sc_hd__buf_6 fanout1385 (.A(net39),
    .X(net1385));
 sky130_fd_sc_hd__buf_2 fanout1418 (.A(net1419),
    .X(net1418));
 sky130_fd_sc_hd__buf_2 fanout1419 (.A(net1420),
    .X(net1419));
 sky130_fd_sc_hd__clkbuf_4 fanout1420 (.A(net1422),
    .X(net1420));
 sky130_fd_sc_hd__buf_4 fanout1421 (.A(net1422),
    .X(net1421));
 sky130_fd_sc_hd__buf_4 fanout1422 (.A(net129),
    .X(net1422));
 sky130_fd_sc_hd__buf_4 fanout1423 (.A(net1424),
    .X(net1423));
 sky130_fd_sc_hd__buf_2 fanout1425 (.A(net1427),
    .X(net1425));
 sky130_fd_sc_hd__clkbuf_2 fanout1426 (.A(net1427),
    .X(net1426));
 sky130_fd_sc_hd__buf_4 fanout1427 (.A(net1430),
    .X(net1427));
 sky130_fd_sc_hd__buf_4 fanout1428 (.A(net1432),
    .X(net1428));
 sky130_fd_sc_hd__buf_4 fanout1429 (.A(net1431),
    .X(net1429));
 sky130_fd_sc_hd__clkbuf_1 fanout1430 (.A(net128),
    .X(net1430));
 sky130_fd_sc_hd__clkbuf_4 fanout1433 (.A(net1435),
    .X(net1433));
 sky130_fd_sc_hd__clkbuf_2 fanout1434 (.A(net1435),
    .X(net1434));
 sky130_fd_sc_hd__buf_4 fanout1435 (.A(net1440),
    .X(net1435));
 sky130_fd_sc_hd__clkbuf_4 fanout1436 (.A(net1440),
    .X(net1436));
 sky130_fd_sc_hd__buf_6 fanout1437 (.A(net1438),
    .X(net1437));
 sky130_fd_sc_hd__buf_6 fanout1438 (.A(net1440),
    .X(net1438));
 sky130_fd_sc_hd__buf_4 fanout1440 (.A(net127),
    .X(net1440));
 sky130_fd_sc_hd__clkbuf_4 fanout1441 (.A(net1443),
    .X(net1441));
 sky130_fd_sc_hd__clkbuf_2 fanout1442 (.A(net1443),
    .X(net1442));
 sky130_fd_sc_hd__buf_4 fanout1443 (.A(net1445),
    .X(net1443));
 sky130_fd_sc_hd__clkbuf_4 fanout1444 (.A(net1445),
    .X(net1444));
 sky130_fd_sc_hd__buf_4 fanout1445 (.A(net126),
    .X(net1445));
 sky130_fd_sc_hd__buf_6 fanout1446 (.A(net1447),
    .X(net1446));
 sky130_fd_sc_hd__buf_6 fanout1447 (.A(net126),
    .X(net1447));
 sky130_fd_sc_hd__clkbuf_4 fanout1448 (.A(net1452),
    .X(net1448));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1449 (.A(net1452),
    .X(net1449));
 sky130_fd_sc_hd__clkbuf_4 fanout1450 (.A(net1451),
    .X(net1450));
 sky130_fd_sc_hd__buf_4 fanout1451 (.A(net1452),
    .X(net1451));
 sky130_fd_sc_hd__clkbuf_4 fanout1452 (.A(net1456),
    .X(net1452));
 sky130_fd_sc_hd__buf_4 fanout1453 (.A(net1455),
    .X(net1453));
 sky130_fd_sc_hd__buf_6 fanout1454 (.A(net1456),
    .X(net1454));
 sky130_fd_sc_hd__clkbuf_4 fanout1457 (.A(net1458),
    .X(net1457));
 sky130_fd_sc_hd__buf_2 fanout1458 (.A(net1459),
    .X(net1458));
 sky130_fd_sc_hd__buf_4 fanout1459 (.A(net1465),
    .X(net1459));
 sky130_fd_sc_hd__clkbuf_4 fanout1460 (.A(net1461),
    .X(net1460));
 sky130_fd_sc_hd__buf_4 fanout1461 (.A(net1465),
    .X(net1461));
 sky130_fd_sc_hd__buf_4 fanout1462 (.A(net1463),
    .X(net1462));
 sky130_fd_sc_hd__clkbuf_1 fanout1463 (.A(net1465),
    .X(net1463));
 sky130_fd_sc_hd__clkbuf_4 fanout1466 (.A(net1467),
    .X(net1466));
 sky130_fd_sc_hd__buf_4 fanout1467 (.A(net1469),
    .X(net1467));
 sky130_fd_sc_hd__buf_6 fanout1468 (.A(net1469),
    .X(net1468));
 sky130_fd_sc_hd__buf_4 fanout1469 (.A(net1473),
    .X(net1469));
 sky130_fd_sc_hd__buf_4 fanout1470 (.A(net1471),
    .X(net1470));
 sky130_fd_sc_hd__buf_6 fanout1471 (.A(net1473),
    .X(net1471));
 sky130_fd_sc_hd__buf_4 fanout1474 (.A(net1477),
    .X(net1474));
 sky130_fd_sc_hd__clkbuf_2 fanout1475 (.A(net1477),
    .X(net1475));
 sky130_fd_sc_hd__clkbuf_4 fanout1476 (.A(net1477),
    .X(net1476));
 sky130_fd_sc_hd__clkbuf_4 fanout1477 (.A(net1478),
    .X(net1477));
 sky130_fd_sc_hd__buf_4 fanout1478 (.A(net1479),
    .X(net1478));
 sky130_fd_sc_hd__buf_6 fanout1479 (.A(net122),
    .X(net1479));
 sky130_fd_sc_hd__clkbuf_4 fanout1481 (.A(net1485),
    .X(net1481));
 sky130_fd_sc_hd__clkbuf_2 fanout1482 (.A(net1485),
    .X(net1482));
 sky130_fd_sc_hd__clkbuf_4 fanout1483 (.A(net1485),
    .X(net1483));
 sky130_fd_sc_hd__clkbuf_4 fanout1484 (.A(net1485),
    .X(net1484));
 sky130_fd_sc_hd__clkbuf_4 fanout1485 (.A(net1486),
    .X(net1485));
 sky130_fd_sc_hd__buf_6 fanout1486 (.A(net121),
    .X(net1486));
 sky130_fd_sc_hd__clkbuf_4 fanout1488 (.A(net1489),
    .X(net1488));
 sky130_fd_sc_hd__clkbuf_2 fanout1489 (.A(net1496),
    .X(net1489));
 sky130_fd_sc_hd__buf_2 fanout1490 (.A(net1492),
    .X(net1490));
 sky130_fd_sc_hd__clkbuf_2 fanout1491 (.A(net1492),
    .X(net1491));
 sky130_fd_sc_hd__buf_4 fanout1492 (.A(net1496),
    .X(net1492));
 sky130_fd_sc_hd__buf_4 fanout1493 (.A(net1494),
    .X(net1493));
 sky130_fd_sc_hd__buf_6 fanout1494 (.A(net1496),
    .X(net1494));
 sky130_fd_sc_hd__buf_4 fanout1496 (.A(net120),
    .X(net1496));
 sky130_fd_sc_hd__buf_2 fanout1498 (.A(net1499),
    .X(net1498));
 sky130_fd_sc_hd__buf_4 fanout1499 (.A(net1502),
    .X(net1499));
 sky130_fd_sc_hd__clkbuf_4 fanout1500 (.A(net1501),
    .X(net1500));
 sky130_fd_sc_hd__clkbuf_4 fanout1501 (.A(net1502),
    .X(net1501));
 sky130_fd_sc_hd__clkbuf_4 fanout1502 (.A(net1503),
    .X(net1502));
 sky130_fd_sc_hd__buf_6 fanout1503 (.A(net119),
    .X(net1503));
 sky130_fd_sc_hd__clkbuf_4 fanout1505 (.A(net1507),
    .X(net1505));
 sky130_fd_sc_hd__clkbuf_2 fanout1506 (.A(net1507),
    .X(net1506));
 sky130_fd_sc_hd__buf_4 fanout1507 (.A(net1509),
    .X(net1507));
 sky130_fd_sc_hd__clkbuf_4 fanout1508 (.A(net1509),
    .X(net1508));
 sky130_fd_sc_hd__buf_4 fanout1509 (.A(net1510),
    .X(net1509));
 sky130_fd_sc_hd__buf_6 fanout1510 (.A(net118),
    .X(net1510));
 sky130_fd_sc_hd__buf_4 fanout1512 (.A(net1515),
    .X(net1512));
 sky130_fd_sc_hd__buf_2 fanout1513 (.A(net1515),
    .X(net1513));
 sky130_fd_sc_hd__clkbuf_4 fanout1514 (.A(net1515),
    .X(net1514));
 sky130_fd_sc_hd__clkbuf_4 fanout1515 (.A(net1516),
    .X(net1515));
 sky130_fd_sc_hd__buf_4 fanout1516 (.A(net1517),
    .X(net1516));
 sky130_fd_sc_hd__buf_6 fanout1517 (.A(net117),
    .X(net1517));
 sky130_fd_sc_hd__buf_2 fanout1519 (.A(net1522),
    .X(net1519));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout1520 (.A(net1522),
    .X(net1520));
 sky130_fd_sc_hd__clkbuf_4 fanout1521 (.A(net1522),
    .X(net1521));
 sky130_fd_sc_hd__buf_4 fanout1522 (.A(net1523),
    .X(net1522));
 sky130_fd_sc_hd__buf_4 fanout1523 (.A(net1524),
    .X(net1523));
 sky130_fd_sc_hd__buf_6 fanout1524 (.A(net116),
    .X(net1524));
 sky130_fd_sc_hd__clkbuf_4 fanout1526 (.A(net1529),
    .X(net1526));
 sky130_fd_sc_hd__clkbuf_2 fanout1527 (.A(net1529),
    .X(net1527));
 sky130_fd_sc_hd__clkbuf_4 fanout1528 (.A(net1529),
    .X(net1528));
 sky130_fd_sc_hd__clkbuf_4 fanout1529 (.A(net1530),
    .X(net1529));
 sky130_fd_sc_hd__clkbuf_8 fanout1530 (.A(net1531),
    .X(net1530));
 sky130_fd_sc_hd__clkbuf_2 fanout1531 (.A(net115),
    .X(net1531));
 sky130_fd_sc_hd__clkbuf_4 fanout1534 (.A(net1535),
    .X(net1534));
 sky130_fd_sc_hd__clkbuf_2 fanout1535 (.A(net1537),
    .X(net1535));
 sky130_fd_sc_hd__clkbuf_4 fanout1536 (.A(net1537),
    .X(net1536));
 sky130_fd_sc_hd__buf_2 fanout1537 (.A(net1538),
    .X(net1537));
 sky130_fd_sc_hd__buf_4 fanout1538 (.A(net1539),
    .X(net1538));
 sky130_fd_sc_hd__buf_6 fanout1539 (.A(net114),
    .X(net1539));
 sky130_fd_sc_hd__clkbuf_4 fanout1541 (.A(net1542),
    .X(net1541));
 sky130_fd_sc_hd__buf_4 fanout1542 (.A(net1543),
    .X(net1542));
 sky130_fd_sc_hd__clkbuf_1 fanout1543 (.A(net113),
    .X(net1543));
 sky130_fd_sc_hd__clkbuf_4 fanout1545 (.A(net1547),
    .X(net1545));
 sky130_fd_sc_hd__buf_4 fanout1546 (.A(net1547),
    .X(net1546));
 sky130_fd_sc_hd__buf_6 fanout1547 (.A(net113),
    .X(net1547));
 sky130_fd_sc_hd__clkbuf_4 fanout1549 (.A(net1550),
    .X(net1549));
 sky130_fd_sc_hd__clkbuf_4 fanout1550 (.A(net1555),
    .X(net1550));
 sky130_fd_sc_hd__buf_4 fanout1551 (.A(net1555),
    .X(net1551));
 sky130_fd_sc_hd__clkbuf_1 fanout1552 (.A(net1555),
    .X(net1552));
 sky130_fd_sc_hd__buf_4 fanout1553 (.A(net1554),
    .X(net1553));
 sky130_fd_sc_hd__buf_4 fanout1554 (.A(net1555),
    .X(net1554));
 sky130_fd_sc_hd__buf_6 fanout1555 (.A(net112),
    .X(net1555));
 sky130_fd_sc_hd__buf_4 fanout1556 (.A(net1557),
    .X(net1556));
 sky130_fd_sc_hd__buf_6 fanout1557 (.A(net111),
    .X(net1557));
 sky130_fd_sc_hd__clkbuf_4 fanout1559 (.A(net1560),
    .X(net1559));
 sky130_fd_sc_hd__clkbuf_4 fanout1560 (.A(net1562),
    .X(net1560));
 sky130_fd_sc_hd__clkbuf_4 fanout1561 (.A(net1563),
    .X(net1561));
 sky130_fd_sc_hd__clkbuf_1 fanout1562 (.A(net111),
    .X(net1562));
 sky130_fd_sc_hd__buf_6 fanout1564 (.A(net110),
    .X(net1564));
 sky130_fd_sc_hd__buf_2 fanout1565 (.A(net110),
    .X(net1565));
 sky130_fd_sc_hd__clkbuf_4 fanout1566 (.A(net1569),
    .X(net1566));
 sky130_fd_sc_hd__clkbuf_2 fanout1567 (.A(net1569),
    .X(net1567));
 sky130_fd_sc_hd__clkbuf_4 fanout1568 (.A(net1569),
    .X(net1568));
 sky130_fd_sc_hd__buf_6 fanout1569 (.A(net110),
    .X(net1569));
 sky130_fd_sc_hd__buf_4 fanout1572 (.A(net1573),
    .X(net1572));
 sky130_fd_sc_hd__buf_4 fanout1573 (.A(net109),
    .X(net1573));
 sky130_fd_sc_hd__buf_4 fanout1574 (.A(net1575),
    .X(net1574));
 sky130_fd_sc_hd__buf_4 fanout1575 (.A(net109),
    .X(net1575));
 sky130_fd_sc_hd__buf_6 fanout1576 (.A(net1577),
    .X(net1576));
 sky130_fd_sc_hd__buf_6 fanout1577 (.A(net109),
    .X(net1577));
 sky130_fd_sc_hd__buf_4 fanout1579 (.A(net108),
    .X(net1579));
 sky130_fd_sc_hd__buf_2 fanout1580 (.A(net108),
    .X(net1580));
 sky130_fd_sc_hd__buf_2 fanout1581 (.A(net1582),
    .X(net1581));
 sky130_fd_sc_hd__clkbuf_4 fanout1582 (.A(net1584),
    .X(net1582));
 sky130_fd_sc_hd__buf_4 fanout1583 (.A(net1585),
    .X(net1583));
 sky130_fd_sc_hd__clkbuf_1 fanout1584 (.A(net108),
    .X(net1584));
 sky130_fd_sc_hd__buf_4 fanout1586 (.A(net1587),
    .X(net1586));
 sky130_fd_sc_hd__buf_6 fanout1587 (.A(net107),
    .X(net1587));
 sky130_fd_sc_hd__clkbuf_4 fanout1589 (.A(net1592),
    .X(net1589));
 sky130_fd_sc_hd__clkbuf_2 fanout1590 (.A(net1592),
    .X(net1590));
 sky130_fd_sc_hd__clkbuf_8 fanout1591 (.A(net1593),
    .X(net1591));
 sky130_fd_sc_hd__buf_6 fanout1592 (.A(net107),
    .X(net1592));
 sky130_fd_sc_hd__buf_6 fanout1595 (.A(net1602),
    .X(net1595));
 sky130_fd_sc_hd__buf_2 fanout1597 (.A(net1602),
    .X(net1597));
 sky130_fd_sc_hd__buf_4 fanout1598 (.A(net1602),
    .X(net1598));
 sky130_fd_sc_hd__clkbuf_2 fanout1599 (.A(net1602),
    .X(net1599));
 sky130_fd_sc_hd__clkbuf_4 fanout1600 (.A(net1601),
    .X(net1600));
 sky130_fd_sc_hd__buf_4 fanout1601 (.A(net1602),
    .X(net1601));
 sky130_fd_sc_hd__buf_8 fanout1602 (.A(net106),
    .X(net1602));
 sky130_fd_sc_hd__buf_4 fanout1603 (.A(net1604),
    .X(net1603));
 sky130_fd_sc_hd__buf_6 fanout1604 (.A(net1610),
    .X(net1604));
 sky130_fd_sc_hd__buf_4 fanout1606 (.A(net1611),
    .X(net1606));
 sky130_fd_sc_hd__buf_4 fanout1607 (.A(net1608),
    .X(net1607));
 sky130_fd_sc_hd__clkbuf_1 fanout1608 (.A(net1611),
    .X(net1608));
 sky130_fd_sc_hd__buf_6 fanout1610 (.A(net105),
    .X(net1610));
 sky130_fd_sc_hd__buf_6 fanout1613 (.A(net1617),
    .X(net1613));
 sky130_fd_sc_hd__buf_2 fanout1614 (.A(net1616),
    .X(net1614));
 sky130_fd_sc_hd__buf_2 fanout1615 (.A(net1616),
    .X(net1615));
 sky130_fd_sc_hd__buf_4 fanout1616 (.A(net1617),
    .X(net1616));
 sky130_fd_sc_hd__buf_4 fanout1617 (.A(net1619),
    .X(net1617));
 sky130_fd_sc_hd__buf_6 fanout1618 (.A(net1620),
    .X(net1618));
 sky130_fd_sc_hd__buf_6 fanout1619 (.A(net104),
    .X(net1619));
 sky130_fd_sc_hd__clkbuf_4 fanout1621 (.A(net1626),
    .X(net1621));
 sky130_fd_sc_hd__clkbuf_2 fanout1622 (.A(net1623),
    .X(net1622));
 sky130_fd_sc_hd__buf_4 fanout1623 (.A(net1626),
    .X(net1623));
 sky130_fd_sc_hd__buf_4 fanout1624 (.A(net1626),
    .X(net1624));
 sky130_fd_sc_hd__buf_4 fanout1625 (.A(net1627),
    .X(net1625));
 sky130_fd_sc_hd__buf_6 fanout1626 (.A(net103),
    .X(net1626));
 sky130_fd_sc_hd__buf_2 fanout1628 (.A(net1630),
    .X(net1628));
 sky130_fd_sc_hd__clkbuf_2 fanout1629 (.A(net1630),
    .X(net1629));
 sky130_fd_sc_hd__buf_4 fanout1630 (.A(net1633),
    .X(net1630));
 sky130_fd_sc_hd__buf_4 fanout1631 (.A(net1635),
    .X(net1631));
 sky130_fd_sc_hd__buf_4 fanout1632 (.A(net1634),
    .X(net1632));
 sky130_fd_sc_hd__clkbuf_1 fanout1633 (.A(net102),
    .X(net1633));
 sky130_fd_sc_hd__clkbuf_4 fanout1636 (.A(net1641),
    .X(net1636));
 sky130_fd_sc_hd__clkbuf_2 fanout1637 (.A(net1638),
    .X(net1637));
 sky130_fd_sc_hd__clkbuf_4 fanout1638 (.A(net1641),
    .X(net1638));
 sky130_fd_sc_hd__buf_4 fanout1639 (.A(net1641),
    .X(net1639));
 sky130_fd_sc_hd__buf_4 fanout1640 (.A(net1642),
    .X(net1640));
 sky130_fd_sc_hd__buf_6 fanout1641 (.A(net101),
    .X(net1641));
 sky130_fd_sc_hd__buf_2 fanout1643 (.A(net1644),
    .X(net1643));
 sky130_fd_sc_hd__buf_4 fanout1644 (.A(net1645),
    .X(net1644));
 sky130_fd_sc_hd__clkbuf_2 fanout1645 (.A(net1648),
    .X(net1645));
 sky130_fd_sc_hd__buf_4 fanout1646 (.A(net1648),
    .X(net1646));
 sky130_fd_sc_hd__buf_4 fanout1647 (.A(net1649),
    .X(net1647));
 sky130_fd_sc_hd__buf_6 fanout1648 (.A(net100),
    .X(net1648));
 sky130_fd_sc_hd__buf_6 fanout1651 (.A(net1),
    .X(net1651));
 sky130_fd_sc_hd__buf_2 fanout513 (.A(_04006_),
    .X(net513));
 sky130_fd_sc_hd__clkbuf_1 fanout514 (.A(_04006_),
    .X(net514));
 sky130_fd_sc_hd__clkbuf_4 fanout515 (.A(_01355_),
    .X(net515));
 sky130_fd_sc_hd__buf_2 fanout516 (.A(_01355_),
    .X(net516));
 sky130_fd_sc_hd__clkbuf_2 fanout517 (.A(net518),
    .X(net517));
 sky130_fd_sc_hd__clkbuf_2 fanout518 (.A(_04039_),
    .X(net518));
 sky130_fd_sc_hd__clkbuf_4 fanout519 (.A(_01348_),
    .X(net519));
 sky130_fd_sc_hd__buf_2 fanout520 (.A(_01348_),
    .X(net520));
 sky130_fd_sc_hd__clkbuf_4 fanout521 (.A(_01343_),
    .X(net521));
 sky130_fd_sc_hd__buf_2 fanout522 (.A(_01343_),
    .X(net522));
 sky130_fd_sc_hd__clkbuf_2 fanout523 (.A(_04072_),
    .X(net523));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout524 (.A(_04072_),
    .X(net524));
 sky130_fd_sc_hd__buf_2 fanout525 (.A(_03763_),
    .X(net525));
 sky130_fd_sc_hd__buf_2 fanout526 (.A(_03703_),
    .X(net526));
 sky130_fd_sc_hd__clkbuf_8 fanout534 (.A(_01032_),
    .X(net534));
 sky130_fd_sc_hd__buf_2 fanout535 (.A(_01032_),
    .X(net535));
 sky130_fd_sc_hd__clkbuf_4 fanout539 (.A(_03524_),
    .X(net539));
 sky130_fd_sc_hd__clkbuf_4 fanout540 (.A(_03524_),
    .X(net540));
 sky130_fd_sc_hd__buf_4 fanout541 (.A(net545),
    .X(net541));
 sky130_fd_sc_hd__buf_2 fanout542 (.A(net544),
    .X(net542));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout543 (.A(net544),
    .X(net543));
 sky130_fd_sc_hd__buf_2 fanout544 (.A(net545),
    .X(net544));
 sky130_fd_sc_hd__buf_2 fanout545 (.A(_03477_),
    .X(net545));
 sky130_fd_sc_hd__clkbuf_4 fanout546 (.A(net547),
    .X(net546));
 sky130_fd_sc_hd__clkbuf_4 fanout547 (.A(_03475_),
    .X(net547));
 sky130_fd_sc_hd__clkbuf_4 fanout548 (.A(_03475_),
    .X(net548));
 sky130_fd_sc_hd__buf_2 fanout549 (.A(_03472_),
    .X(net549));
 sky130_fd_sc_hd__clkbuf_1 fanout550 (.A(_03472_),
    .X(net550));
 sky130_fd_sc_hd__buf_2 fanout551 (.A(net552),
    .X(net551));
 sky130_fd_sc_hd__clkbuf_2 fanout552 (.A(_03471_),
    .X(net552));
 sky130_fd_sc_hd__clkbuf_4 fanout553 (.A(_03470_),
    .X(net553));
 sky130_fd_sc_hd__clkbuf_2 fanout554 (.A(_03470_),
    .X(net554));
 sky130_fd_sc_hd__buf_2 fanout555 (.A(_03470_),
    .X(net555));
 sky130_fd_sc_hd__buf_2 fanout556 (.A(_03470_),
    .X(net556));
 sky130_fd_sc_hd__buf_2 fanout557 (.A(net558),
    .X(net557));
 sky130_fd_sc_hd__buf_2 fanout558 (.A(_03466_),
    .X(net558));
 sky130_fd_sc_hd__buf_2 fanout559 (.A(_03464_),
    .X(net559));
 sky130_fd_sc_hd__clkbuf_4 fanout560 (.A(net561),
    .X(net560));
 sky130_fd_sc_hd__buf_4 fanout561 (.A(net563),
    .X(net561));
 sky130_fd_sc_hd__clkbuf_4 fanout562 (.A(net563),
    .X(net562));
 sky130_fd_sc_hd__clkbuf_4 fanout563 (.A(_01785_),
    .X(net563));
 sky130_fd_sc_hd__clkbuf_4 fanout568 (.A(net569),
    .X(net568));
 sky130_fd_sc_hd__clkbuf_4 fanout569 (.A(_01239_),
    .X(net569));
 sky130_fd_sc_hd__clkbuf_4 fanout570 (.A(_01239_),
    .X(net570));
 sky130_fd_sc_hd__clkbuf_4 fanout571 (.A(net573),
    .X(net571));
 sky130_fd_sc_hd__clkbuf_2 fanout572 (.A(net573),
    .X(net572));
 sky130_fd_sc_hd__buf_2 fanout573 (.A(net574),
    .X(net573));
 sky130_fd_sc_hd__clkbuf_4 fanout574 (.A(_01198_),
    .X(net574));
 sky130_fd_sc_hd__buf_4 fanout575 (.A(_01005_),
    .X(net575));
 sky130_fd_sc_hd__buf_2 fanout576 (.A(_01005_),
    .X(net576));
 sky130_fd_sc_hd__buf_4 fanout577 (.A(net578),
    .X(net577));
 sky130_fd_sc_hd__buf_4 fanout578 (.A(_01005_),
    .X(net578));
 sky130_fd_sc_hd__clkbuf_4 fanout579 (.A(_04312_),
    .X(net579));
 sky130_fd_sc_hd__clkbuf_2 fanout580 (.A(_04312_),
    .X(net580));
 sky130_fd_sc_hd__buf_2 fanout584 (.A(net586),
    .X(net584));
 sky130_fd_sc_hd__clkbuf_2 fanout585 (.A(net586),
    .X(net585));
 sky130_fd_sc_hd__clkbuf_4 fanout586 (.A(_03478_),
    .X(net586));
 sky130_fd_sc_hd__buf_2 fanout587 (.A(_03041_),
    .X(net587));
 sky130_fd_sc_hd__buf_2 fanout588 (.A(_03038_),
    .X(net588));
 sky130_fd_sc_hd__buf_4 fanout589 (.A(net590),
    .X(net589));
 sky130_fd_sc_hd__clkbuf_4 fanout590 (.A(_01793_),
    .X(net590));
 sky130_fd_sc_hd__clkbuf_4 fanout591 (.A(_01793_),
    .X(net591));
 sky130_fd_sc_hd__clkbuf_2 fanout592 (.A(_01793_),
    .X(net592));
 sky130_fd_sc_hd__clkbuf_4 fanout593 (.A(net594),
    .X(net593));
 sky130_fd_sc_hd__clkbuf_4 fanout594 (.A(net595),
    .X(net594));
 sky130_fd_sc_hd__buf_4 fanout595 (.A(_01788_),
    .X(net595));
 sky130_fd_sc_hd__clkbuf_8 fanout596 (.A(_01782_),
    .X(net596));
 sky130_fd_sc_hd__clkbuf_4 fanout597 (.A(_01782_),
    .X(net597));
 sky130_fd_sc_hd__buf_2 fanout598 (.A(net599),
    .X(net598));
 sky130_fd_sc_hd__clkbuf_4 fanout599 (.A(net600),
    .X(net599));
 sky130_fd_sc_hd__buf_2 fanout600 (.A(_01649_),
    .X(net600));
 sky130_fd_sc_hd__buf_4 fanout603 (.A(net604),
    .X(net603));
 sky130_fd_sc_hd__buf_4 fanout604 (.A(net606),
    .X(net604));
 sky130_fd_sc_hd__buf_6 fanout605 (.A(net606),
    .X(net605));
 sky130_fd_sc_hd__buf_6 fanout606 (.A(_01558_),
    .X(net606));
 sky130_fd_sc_hd__buf_4 fanout607 (.A(net609),
    .X(net607));
 sky130_fd_sc_hd__clkbuf_2 fanout608 (.A(net609),
    .X(net608));
 sky130_fd_sc_hd__buf_2 fanout609 (.A(_01557_),
    .X(net609));
 sky130_fd_sc_hd__clkbuf_4 fanout610 (.A(_01557_),
    .X(net610));
 sky130_fd_sc_hd__buf_2 fanout611 (.A(_01557_),
    .X(net611));
 sky130_fd_sc_hd__clkbuf_4 fanout612 (.A(net613),
    .X(net612));
 sky130_fd_sc_hd__buf_4 fanout613 (.A(net615),
    .X(net613));
 sky130_fd_sc_hd__clkbuf_4 fanout614 (.A(net615),
    .X(net614));
 sky130_fd_sc_hd__buf_4 fanout615 (.A(_01556_),
    .X(net615));
 sky130_fd_sc_hd__clkbuf_4 fanout616 (.A(net617),
    .X(net616));
 sky130_fd_sc_hd__clkbuf_4 fanout617 (.A(net619),
    .X(net617));
 sky130_fd_sc_hd__buf_4 fanout618 (.A(net619),
    .X(net618));
 sky130_fd_sc_hd__buf_4 fanout619 (.A(_01555_),
    .X(net619));
 sky130_fd_sc_hd__clkbuf_4 fanout620 (.A(net622),
    .X(net620));
 sky130_fd_sc_hd__clkbuf_4 fanout621 (.A(net622),
    .X(net621));
 sky130_fd_sc_hd__clkbuf_4 fanout622 (.A(_01554_),
    .X(net622));
 sky130_fd_sc_hd__buf_4 fanout623 (.A(_01554_),
    .X(net623));
 sky130_fd_sc_hd__buf_4 fanout624 (.A(_01553_),
    .X(net624));
 sky130_fd_sc_hd__clkbuf_2 fanout625 (.A(_01553_),
    .X(net625));
 sky130_fd_sc_hd__clkbuf_4 fanout626 (.A(net627),
    .X(net626));
 sky130_fd_sc_hd__buf_4 fanout627 (.A(_01553_),
    .X(net627));
 sky130_fd_sc_hd__buf_4 fanout628 (.A(net629),
    .X(net628));
 sky130_fd_sc_hd__buf_4 fanout629 (.A(net632),
    .X(net629));
 sky130_fd_sc_hd__buf_4 fanout630 (.A(net632),
    .X(net630));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout631 (.A(net632),
    .X(net631));
 sky130_fd_sc_hd__clkbuf_4 fanout632 (.A(_01552_),
    .X(net632));
 sky130_fd_sc_hd__clkbuf_4 fanout633 (.A(net634),
    .X(net633));
 sky130_fd_sc_hd__clkbuf_4 fanout634 (.A(_01551_),
    .X(net634));
 sky130_fd_sc_hd__clkbuf_4 fanout635 (.A(net636),
    .X(net635));
 sky130_fd_sc_hd__clkbuf_4 fanout636 (.A(_01551_),
    .X(net636));
 sky130_fd_sc_hd__clkbuf_4 fanout637 (.A(net638),
    .X(net637));
 sky130_fd_sc_hd__buf_4 fanout638 (.A(_01550_),
    .X(net638));
 sky130_fd_sc_hd__clkbuf_4 fanout639 (.A(_01550_),
    .X(net639));
 sky130_fd_sc_hd__clkbuf_2 fanout640 (.A(_01550_),
    .X(net640));
 sky130_fd_sc_hd__buf_4 fanout641 (.A(net642),
    .X(net641));
 sky130_fd_sc_hd__buf_4 fanout642 (.A(net644),
    .X(net642));
 sky130_fd_sc_hd__buf_4 fanout643 (.A(net644),
    .X(net643));
 sky130_fd_sc_hd__buf_4 fanout644 (.A(_01549_),
    .X(net644));
 sky130_fd_sc_hd__clkbuf_4 fanout645 (.A(_01548_),
    .X(net645));
 sky130_fd_sc_hd__clkbuf_4 fanout646 (.A(_01548_),
    .X(net646));
 sky130_fd_sc_hd__clkbuf_4 fanout647 (.A(net648),
    .X(net647));
 sky130_fd_sc_hd__buf_4 fanout648 (.A(_01548_),
    .X(net648));
 sky130_fd_sc_hd__buf_4 fanout649 (.A(net651),
    .X(net649));
 sky130_fd_sc_hd__buf_2 fanout650 (.A(net651),
    .X(net650));
 sky130_fd_sc_hd__clkbuf_4 fanout651 (.A(net653),
    .X(net651));
 sky130_fd_sc_hd__buf_4 fanout652 (.A(net653),
    .X(net652));
 sky130_fd_sc_hd__clkbuf_4 fanout653 (.A(_01547_),
    .X(net653));
 sky130_fd_sc_hd__clkbuf_4 fanout654 (.A(net656),
    .X(net654));
 sky130_fd_sc_hd__buf_2 fanout655 (.A(net656),
    .X(net655));
 sky130_fd_sc_hd__clkbuf_4 fanout656 (.A(net658),
    .X(net656));
 sky130_fd_sc_hd__buf_4 fanout657 (.A(net658),
    .X(net657));
 sky130_fd_sc_hd__clkbuf_4 fanout658 (.A(_01545_),
    .X(net658));
 sky130_fd_sc_hd__buf_4 fanout659 (.A(net660),
    .X(net659));
 sky130_fd_sc_hd__buf_4 fanout660 (.A(net663),
    .X(net660));
 sky130_fd_sc_hd__buf_4 fanout661 (.A(net663),
    .X(net661));
 sky130_fd_sc_hd__buf_2 fanout662 (.A(net663),
    .X(net662));
 sky130_fd_sc_hd__buf_4 fanout663 (.A(_01542_),
    .X(net663));
 sky130_fd_sc_hd__buf_4 fanout664 (.A(net665),
    .X(net664));
 sky130_fd_sc_hd__buf_4 fanout665 (.A(_01539_),
    .X(net665));
 sky130_fd_sc_hd__clkbuf_4 fanout666 (.A(net667),
    .X(net666));
 sky130_fd_sc_hd__clkbuf_4 fanout667 (.A(_01539_),
    .X(net667));
 sky130_fd_sc_hd__buf_4 fanout668 (.A(net669),
    .X(net668));
 sky130_fd_sc_hd__clkbuf_4 fanout669 (.A(_01538_),
    .X(net669));
 sky130_fd_sc_hd__buf_6 fanout670 (.A(_01538_),
    .X(net670));
 sky130_fd_sc_hd__buf_2 fanout671 (.A(_01538_),
    .X(net671));
 sky130_fd_sc_hd__buf_2 fanout672 (.A(net673),
    .X(net672));
 sky130_fd_sc_hd__clkbuf_2 fanout673 (.A(_01501_),
    .X(net673));
 sky130_fd_sc_hd__buf_2 fanout674 (.A(_01482_),
    .X(net674));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout675 (.A(_01482_),
    .X(net675));
 sky130_fd_sc_hd__clkbuf_2 fanout676 (.A(_01463_),
    .X(net676));
 sky130_fd_sc_hd__clkbuf_2 fanout677 (.A(_01463_),
    .X(net677));
 sky130_fd_sc_hd__clkbuf_4 fanout678 (.A(net680),
    .X(net678));
 sky130_fd_sc_hd__clkbuf_2 fanout679 (.A(net680),
    .X(net679));
 sky130_fd_sc_hd__buf_2 fanout680 (.A(_01334_),
    .X(net680));
 sky130_fd_sc_hd__buf_2 fanout681 (.A(net683),
    .X(net681));
 sky130_fd_sc_hd__clkbuf_2 fanout682 (.A(net683),
    .X(net682));
 sky130_fd_sc_hd__buf_4 fanout683 (.A(_01146_),
    .X(net683));
 sky130_fd_sc_hd__clkbuf_4 fanout684 (.A(_01146_),
    .X(net684));
 sky130_fd_sc_hd__clkbuf_4 fanout685 (.A(net690),
    .X(net685));
 sky130_fd_sc_hd__clkbuf_2 fanout686 (.A(net690),
    .X(net686));
 sky130_fd_sc_hd__clkbuf_4 fanout687 (.A(net688),
    .X(net687));
 sky130_fd_sc_hd__clkbuf_2 fanout688 (.A(net689),
    .X(net688));
 sky130_fd_sc_hd__buf_2 fanout689 (.A(net690),
    .X(net689));
 sky130_fd_sc_hd__clkbuf_4 fanout690 (.A(_01134_),
    .X(net690));
 sky130_fd_sc_hd__clkbuf_4 fanout691 (.A(net692),
    .X(net691));
 sky130_fd_sc_hd__buf_2 fanout692 (.A(net693),
    .X(net692));
 sky130_fd_sc_hd__buf_4 fanout693 (.A(_01133_),
    .X(net693));
 sky130_fd_sc_hd__buf_2 fanout694 (.A(net695),
    .X(net694));
 sky130_fd_sc_hd__clkbuf_4 fanout695 (.A(net696),
    .X(net695));
 sky130_fd_sc_hd__clkbuf_4 fanout696 (.A(net697),
    .X(net696));
 sky130_fd_sc_hd__buf_4 fanout697 (.A(_01133_),
    .X(net697));
 sky130_fd_sc_hd__buf_4 fanout698 (.A(_01132_),
    .X(net698));
 sky130_fd_sc_hd__clkbuf_4 fanout699 (.A(_01132_),
    .X(net699));
 sky130_fd_sc_hd__clkbuf_4 fanout700 (.A(_01132_),
    .X(net700));
 sky130_fd_sc_hd__clkbuf_4 fanout701 (.A(_01132_),
    .X(net701));
 sky130_fd_sc_hd__clkbuf_4 fanout702 (.A(net703),
    .X(net702));
 sky130_fd_sc_hd__buf_4 fanout703 (.A(net704),
    .X(net703));
 sky130_fd_sc_hd__buf_4 fanout704 (.A(_01131_),
    .X(net704));
 sky130_fd_sc_hd__clkbuf_4 fanout705 (.A(net706),
    .X(net705));
 sky130_fd_sc_hd__buf_2 fanout706 (.A(net707),
    .X(net706));
 sky130_fd_sc_hd__buf_6 fanout707 (.A(_01131_),
    .X(net707));
 sky130_fd_sc_hd__clkbuf_4 fanout708 (.A(net710),
    .X(net708));
 sky130_fd_sc_hd__buf_2 fanout709 (.A(net710),
    .X(net709));
 sky130_fd_sc_hd__buf_2 fanout710 (.A(net711),
    .X(net710));
 sky130_fd_sc_hd__buf_4 fanout711 (.A(_01008_),
    .X(net711));
 sky130_fd_sc_hd__buf_2 fanout712 (.A(net713),
    .X(net712));
 sky130_fd_sc_hd__buf_2 fanout713 (.A(net714),
    .X(net713));
 sky130_fd_sc_hd__buf_2 fanout714 (.A(_01001_),
    .X(net714));
 sky130_fd_sc_hd__clkbuf_4 fanout715 (.A(_01000_),
    .X(net715));
 sky130_fd_sc_hd__clkbuf_4 fanout716 (.A(_01000_),
    .X(net716));
 sky130_fd_sc_hd__buf_4 fanout717 (.A(_01000_),
    .X(net717));
 sky130_fd_sc_hd__clkbuf_2 fanout718 (.A(_01000_),
    .X(net718));
 sky130_fd_sc_hd__buf_4 fanout719 (.A(net720),
    .X(net719));
 sky130_fd_sc_hd__clkbuf_2 fanout720 (.A(_00250_),
    .X(net720));
 sky130_fd_sc_hd__buf_6 fanout722 (.A(_00250_),
    .X(net722));
 sky130_fd_sc_hd__buf_2 fanout723 (.A(_00985_),
    .X(net723));
 sky130_fd_sc_hd__dlymetal6s2s_1 fanout724 (.A(_00985_),
    .X(net724));
 sky130_fd_sc_hd__buf_2 fanout725 (.A(_00911_),
    .X(net725));
 sky130_fd_sc_hd__clkbuf_4 fanout726 (.A(_00888_),
    .X(net726));
 sky130_fd_sc_hd__buf_2 fanout727 (.A(_00878_),
    .X(net727));
 sky130_fd_sc_hd__buf_2 fanout728 (.A(_00867_),
    .X(net728));
 sky130_fd_sc_hd__clkbuf_4 fanout729 (.A(net730),
    .X(net729));
 sky130_fd_sc_hd__buf_2 fanout730 (.A(_00837_),
    .X(net730));
 sky130_fd_sc_hd__clkbuf_4 fanout731 (.A(_00837_),
    .X(net731));
 sky130_fd_sc_hd__clkbuf_4 fanout732 (.A(net733),
    .X(net732));
 sky130_fd_sc_hd__clkbuf_4 fanout733 (.A(net734),
    .X(net733));
 sky130_fd_sc_hd__clkbuf_4 fanout734 (.A(_00813_),
    .X(net734));
 sky130_fd_sc_hd__buf_2 fanout735 (.A(net738),
    .X(net735));
 sky130_fd_sc_hd__clkbuf_4 fanout736 (.A(net737),
    .X(net736));
 sky130_fd_sc_hd__clkbuf_4 fanout737 (.A(net738),
    .X(net737));
 sky130_fd_sc_hd__buf_2 fanout738 (.A(net751),
    .X(net738));
 sky130_fd_sc_hd__clkbuf_4 fanout739 (.A(net740),
    .X(net739));
 sky130_fd_sc_hd__clkbuf_4 fanout740 (.A(net743),
    .X(net740));
 sky130_fd_sc_hd__clkbuf_4 fanout741 (.A(net742),
    .X(net741));
 sky130_fd_sc_hd__clkbuf_4 fanout742 (.A(net743),
    .X(net742));
 sky130_fd_sc_hd__clkbuf_2 fanout743 (.A(net751),
    .X(net743));
 sky130_fd_sc_hd__buf_4 fanout744 (.A(net746),
    .X(net744));
 sky130_fd_sc_hd__clkbuf_4 fanout745 (.A(net746),
    .X(net745));
 sky130_fd_sc_hd__clkbuf_4 fanout746 (.A(net751),
    .X(net746));
 sky130_fd_sc_hd__clkbuf_4 fanout747 (.A(net748),
    .X(net747));
 sky130_fd_sc_hd__clkbuf_4 fanout748 (.A(net751),
    .X(net748));
 sky130_fd_sc_hd__clkbuf_4 fanout749 (.A(net751),
    .X(net749));
 sky130_fd_sc_hd__clkbuf_2 fanout750 (.A(net751),
    .X(net750));
 sky130_fd_sc_hd__clkbuf_4 fanout751 (.A(net772),
    .X(net751));
 sky130_fd_sc_hd__clkbuf_4 fanout752 (.A(net755),
    .X(net752));
 sky130_fd_sc_hd__clkbuf_4 fanout753 (.A(net754),
    .X(net753));
 sky130_fd_sc_hd__clkbuf_4 fanout754 (.A(net755),
    .X(net754));
 sky130_fd_sc_hd__clkbuf_2 fanout755 (.A(net772),
    .X(net755));
 sky130_fd_sc_hd__clkbuf_4 fanout756 (.A(net758),
    .X(net756));
 sky130_fd_sc_hd__clkbuf_4 fanout757 (.A(net758),
    .X(net757));
 sky130_fd_sc_hd__clkbuf_4 fanout758 (.A(net772),
    .X(net758));
 sky130_fd_sc_hd__clkbuf_4 fanout759 (.A(net762),
    .X(net759));
 sky130_fd_sc_hd__clkbuf_4 fanout760 (.A(net762),
    .X(net760));
 sky130_fd_sc_hd__clkbuf_2 fanout761 (.A(net762),
    .X(net761));
 sky130_fd_sc_hd__clkbuf_2 fanout762 (.A(net772),
    .X(net762));
 sky130_fd_sc_hd__buf_4 fanout763 (.A(net771),
    .X(net763));
 sky130_fd_sc_hd__clkbuf_4 fanout764 (.A(net771),
    .X(net764));
 sky130_fd_sc_hd__clkbuf_4 fanout765 (.A(net771),
    .X(net765));
 sky130_fd_sc_hd__clkbuf_4 fanout766 (.A(net768),
    .X(net766));
 sky130_fd_sc_hd__clkbuf_4 fanout767 (.A(net768),
    .X(net767));
 sky130_fd_sc_hd__buf_2 fanout768 (.A(net771),
    .X(net768));
 sky130_fd_sc_hd__clkbuf_4 fanout769 (.A(net770),
    .X(net769));
 sky130_fd_sc_hd__clkbuf_4 fanout770 (.A(net771),
    .X(net770));
 sky130_fd_sc_hd__clkbuf_4 fanout771 (.A(net772),
    .X(net771));
 sky130_fd_sc_hd__buf_2 fanout772 (.A(net1042),
    .X(net772));
 sky130_fd_sc_hd__clkbuf_4 fanout773 (.A(net774),
    .X(net773));
 sky130_fd_sc_hd__buf_2 fanout774 (.A(net775),
    .X(net774));
 sky130_fd_sc_hd__clkbuf_4 fanout775 (.A(net789),
    .X(net775));
 sky130_fd_sc_hd__clkbuf_4 fanout776 (.A(net779),
    .X(net776));
 sky130_fd_sc_hd__clkbuf_4 fanout777 (.A(net779),
    .X(net777));
 sky130_fd_sc_hd__clkbuf_2 fanout778 (.A(net779),
    .X(net778));
 sky130_fd_sc_hd__clkbuf_2 fanout779 (.A(net789),
    .X(net779));
 sky130_fd_sc_hd__clkbuf_4 fanout780 (.A(net781),
    .X(net780));
 sky130_fd_sc_hd__clkbuf_4 fanout781 (.A(net789),
    .X(net781));
 sky130_fd_sc_hd__clkbuf_4 fanout782 (.A(net783),
    .X(net782));
 sky130_fd_sc_hd__clkbuf_4 fanout783 (.A(net789),
    .X(net783));
 sky130_fd_sc_hd__clkbuf_4 fanout784 (.A(net788),
    .X(net784));
 sky130_fd_sc_hd__clkbuf_4 fanout785 (.A(net788),
    .X(net785));
 sky130_fd_sc_hd__clkbuf_4 fanout786 (.A(net787),
    .X(net786));
 sky130_fd_sc_hd__clkbuf_4 fanout787 (.A(net788),
    .X(net787));
 sky130_fd_sc_hd__clkbuf_2 fanout788 (.A(net789),
    .X(net788));
 sky130_fd_sc_hd__clkbuf_4 fanout789 (.A(net1042),
    .X(net789));
 sky130_fd_sc_hd__clkbuf_4 fanout790 (.A(net791),
    .X(net790));
 sky130_fd_sc_hd__clkbuf_4 fanout791 (.A(net794),
    .X(net791));
 sky130_fd_sc_hd__clkbuf_4 fanout792 (.A(net793),
    .X(net792));
 sky130_fd_sc_hd__clkbuf_4 fanout793 (.A(net794),
    .X(net793));
 sky130_fd_sc_hd__buf_2 fanout794 (.A(net815),
    .X(net794));
 sky130_fd_sc_hd__clkbuf_4 fanout795 (.A(net797),
    .X(net795));
 sky130_fd_sc_hd__clkbuf_4 fanout796 (.A(net797),
    .X(net796));
 sky130_fd_sc_hd__buf_2 fanout797 (.A(net815),
    .X(net797));
 sky130_fd_sc_hd__clkbuf_4 fanout798 (.A(net800),
    .X(net798));
 sky130_fd_sc_hd__clkbuf_4 fanout799 (.A(net800),
    .X(net799));
 sky130_fd_sc_hd__buf_2 fanout800 (.A(net815),
    .X(net800));
 sky130_fd_sc_hd__clkbuf_4 fanout801 (.A(net803),
    .X(net801));
 sky130_fd_sc_hd__clkbuf_4 fanout802 (.A(net803),
    .X(net802));
 sky130_fd_sc_hd__buf_2 fanout803 (.A(net807),
    .X(net803));
 sky130_fd_sc_hd__clkbuf_4 fanout804 (.A(net807),
    .X(net804));
 sky130_fd_sc_hd__clkbuf_4 fanout805 (.A(net807),
    .X(net805));
 sky130_fd_sc_hd__clkbuf_2 fanout806 (.A(net807),
    .X(net806));
 sky130_fd_sc_hd__clkbuf_2 fanout807 (.A(net815),
    .X(net807));
 sky130_fd_sc_hd__clkbuf_4 fanout808 (.A(net810),
    .X(net808));
 sky130_fd_sc_hd__clkbuf_4 fanout809 (.A(net810),
    .X(net809));
 sky130_fd_sc_hd__buf_2 fanout810 (.A(net814),
    .X(net810));
 sky130_fd_sc_hd__clkbuf_4 fanout811 (.A(net814),
    .X(net811));
 sky130_fd_sc_hd__clkbuf_4 fanout812 (.A(net814),
    .X(net812));
 sky130_fd_sc_hd__buf_2 fanout813 (.A(net814),
    .X(net813));
 sky130_fd_sc_hd__clkbuf_2 fanout814 (.A(net815),
    .X(net814));
 sky130_fd_sc_hd__buf_2 fanout815 (.A(net1042),
    .X(net815));
 sky130_fd_sc_hd__buf_4 fanout816 (.A(net836),
    .X(net816));
 sky130_fd_sc_hd__buf_2 fanout817 (.A(net836),
    .X(net817));
 sky130_fd_sc_hd__clkbuf_4 fanout818 (.A(net821),
    .X(net818));
 sky130_fd_sc_hd__clkbuf_4 fanout819 (.A(net821),
    .X(net819));
 sky130_fd_sc_hd__clkbuf_2 fanout820 (.A(net821),
    .X(net820));
 sky130_fd_sc_hd__buf_2 fanout821 (.A(net836),
    .X(net821));
 sky130_fd_sc_hd__clkbuf_4 fanout822 (.A(net825),
    .X(net822));
 sky130_fd_sc_hd__clkbuf_2 fanout823 (.A(net825),
    .X(net823));
 sky130_fd_sc_hd__clkbuf_4 fanout824 (.A(net825),
    .X(net824));
 sky130_fd_sc_hd__clkbuf_2 fanout825 (.A(net836),
    .X(net825));
 sky130_fd_sc_hd__clkbuf_4 fanout826 (.A(net836),
    .X(net826));
 sky130_fd_sc_hd__clkbuf_2 fanout827 (.A(net828),
    .X(net827));
 sky130_fd_sc_hd__clkbuf_4 fanout828 (.A(net836),
    .X(net828));
 sky130_fd_sc_hd__clkbuf_4 fanout829 (.A(net835),
    .X(net829));
 sky130_fd_sc_hd__clkbuf_2 fanout830 (.A(net835),
    .X(net830));
 sky130_fd_sc_hd__clkbuf_4 fanout831 (.A(net835),
    .X(net831));
 sky130_fd_sc_hd__clkbuf_4 fanout832 (.A(net834),
    .X(net832));
 sky130_fd_sc_hd__clkbuf_4 fanout833 (.A(net834),
    .X(net833));
 sky130_fd_sc_hd__buf_2 fanout834 (.A(net835),
    .X(net834));
 sky130_fd_sc_hd__clkbuf_2 fanout835 (.A(net836),
    .X(net835));
 sky130_fd_sc_hd__clkbuf_4 fanout836 (.A(net851),
    .X(net836));
 sky130_fd_sc_hd__clkbuf_4 fanout837 (.A(net838),
    .X(net837));
 sky130_fd_sc_hd__clkbuf_4 fanout838 (.A(net851),
    .X(net838));
 sky130_fd_sc_hd__clkbuf_4 fanout839 (.A(net840),
    .X(net839));
 sky130_fd_sc_hd__clkbuf_4 fanout840 (.A(net842),
    .X(net840));
 sky130_fd_sc_hd__buf_4 fanout841 (.A(net842),
    .X(net841));
 sky130_fd_sc_hd__clkbuf_2 fanout842 (.A(net851),
    .X(net842));
 sky130_fd_sc_hd__clkbuf_4 fanout843 (.A(net846),
    .X(net843));
 sky130_fd_sc_hd__clkbuf_2 fanout844 (.A(net846),
    .X(net844));
 sky130_fd_sc_hd__clkbuf_4 fanout845 (.A(net846),
    .X(net845));
 sky130_fd_sc_hd__buf_2 fanout846 (.A(net850),
    .X(net846));
 sky130_fd_sc_hd__clkbuf_4 fanout847 (.A(net850),
    .X(net847));
 sky130_fd_sc_hd__clkbuf_2 fanout848 (.A(net850),
    .X(net848));
 sky130_fd_sc_hd__clkbuf_4 fanout849 (.A(net850),
    .X(net849));
 sky130_fd_sc_hd__clkbuf_4 fanout850 (.A(net851),
    .X(net850));
 sky130_fd_sc_hd__buf_2 fanout851 (.A(net897),
    .X(net851));
 sky130_fd_sc_hd__clkbuf_4 fanout852 (.A(net855),
    .X(net852));
 sky130_fd_sc_hd__clkbuf_4 fanout853 (.A(net855),
    .X(net853));
 sky130_fd_sc_hd__clkbuf_2 fanout854 (.A(net855),
    .X(net854));
 sky130_fd_sc_hd__clkbuf_2 fanout855 (.A(net858),
    .X(net855));
 sky130_fd_sc_hd__clkbuf_4 fanout856 (.A(net858),
    .X(net856));
 sky130_fd_sc_hd__clkbuf_4 fanout857 (.A(net858),
    .X(net857));
 sky130_fd_sc_hd__buf_2 fanout858 (.A(net897),
    .X(net858));
 sky130_fd_sc_hd__clkbuf_4 fanout859 (.A(net866),
    .X(net859));
 sky130_fd_sc_hd__clkbuf_2 fanout860 (.A(net866),
    .X(net860));
 sky130_fd_sc_hd__clkbuf_4 fanout861 (.A(net866),
    .X(net861));
 sky130_fd_sc_hd__clkbuf_2 fanout862 (.A(net866),
    .X(net862));
 sky130_fd_sc_hd__clkbuf_4 fanout863 (.A(net865),
    .X(net863));
 sky130_fd_sc_hd__clkbuf_4 fanout864 (.A(net865),
    .X(net864));
 sky130_fd_sc_hd__buf_2 fanout865 (.A(net866),
    .X(net865));
 sky130_fd_sc_hd__clkbuf_2 fanout866 (.A(net897),
    .X(net866));
 sky130_fd_sc_hd__clkbuf_4 fanout867 (.A(net868),
    .X(net867));
 sky130_fd_sc_hd__clkbuf_4 fanout868 (.A(net871),
    .X(net868));
 sky130_fd_sc_hd__clkbuf_4 fanout869 (.A(net870),
    .X(net869));
 sky130_fd_sc_hd__clkbuf_4 fanout870 (.A(net871),
    .X(net870));
 sky130_fd_sc_hd__clkbuf_2 fanout871 (.A(net878),
    .X(net871));
 sky130_fd_sc_hd__clkbuf_4 fanout872 (.A(net878),
    .X(net872));
 sky130_fd_sc_hd__clkbuf_2 fanout873 (.A(net878),
    .X(net873));
 sky130_fd_sc_hd__clkbuf_4 fanout874 (.A(net878),
    .X(net874));
 sky130_fd_sc_hd__clkbuf_4 fanout875 (.A(net877),
    .X(net875));
 sky130_fd_sc_hd__clkbuf_4 fanout876 (.A(net877),
    .X(net876));
 sky130_fd_sc_hd__clkbuf_4 fanout877 (.A(net878),
    .X(net877));
 sky130_fd_sc_hd__clkbuf_2 fanout878 (.A(net897),
    .X(net878));
 sky130_fd_sc_hd__buf_4 fanout879 (.A(net882),
    .X(net879));
 sky130_fd_sc_hd__clkbuf_4 fanout880 (.A(net882),
    .X(net880));
 sky130_fd_sc_hd__clkbuf_2 fanout881 (.A(net882),
    .X(net881));
 sky130_fd_sc_hd__buf_2 fanout882 (.A(net896),
    .X(net882));
 sky130_fd_sc_hd__clkbuf_4 fanout883 (.A(net886),
    .X(net883));
 sky130_fd_sc_hd__clkbuf_4 fanout884 (.A(net886),
    .X(net884));
 sky130_fd_sc_hd__clkbuf_2 fanout885 (.A(net886),
    .X(net885));
 sky130_fd_sc_hd__buf_2 fanout886 (.A(net896),
    .X(net886));
 sky130_fd_sc_hd__clkbuf_4 fanout887 (.A(net889),
    .X(net887));
 sky130_fd_sc_hd__clkbuf_2 fanout888 (.A(net889),
    .X(net888));
 sky130_fd_sc_hd__clkbuf_4 fanout889 (.A(net896),
    .X(net889));
 sky130_fd_sc_hd__clkbuf_4 fanout890 (.A(net891),
    .X(net890));
 sky130_fd_sc_hd__clkbuf_4 fanout891 (.A(net892),
    .X(net891));
 sky130_fd_sc_hd__clkbuf_4 fanout892 (.A(net896),
    .X(net892));
 sky130_fd_sc_hd__clkbuf_4 fanout893 (.A(net895),
    .X(net893));
 sky130_fd_sc_hd__clkbuf_4 fanout894 (.A(net895),
    .X(net894));
 sky130_fd_sc_hd__buf_2 fanout895 (.A(net896),
    .X(net895));
 sky130_fd_sc_hd__buf_2 fanout896 (.A(net897),
    .X(net896));
 sky130_fd_sc_hd__clkbuf_4 fanout897 (.A(net1042),
    .X(net897));
 sky130_fd_sc_hd__buf_4 fanout898 (.A(net901),
    .X(net898));
 sky130_fd_sc_hd__clkbuf_4 fanout899 (.A(net900),
    .X(net899));
 sky130_fd_sc_hd__clkbuf_4 fanout900 (.A(net901),
    .X(net900));
 sky130_fd_sc_hd__clkbuf_4 fanout901 (.A(net906),
    .X(net901));
 sky130_fd_sc_hd__buf_4 fanout902 (.A(net906),
    .X(net902));
 sky130_fd_sc_hd__clkbuf_4 fanout903 (.A(net905),
    .X(net903));
 sky130_fd_sc_hd__clkbuf_4 fanout904 (.A(net905),
    .X(net904));
 sky130_fd_sc_hd__buf_2 fanout905 (.A(net906),
    .X(net905));
 sky130_fd_sc_hd__clkbuf_2 fanout906 (.A(net936),
    .X(net906));
 sky130_fd_sc_hd__clkbuf_4 fanout907 (.A(net908),
    .X(net907));
 sky130_fd_sc_hd__clkbuf_4 fanout908 (.A(net909),
    .X(net908));
 sky130_fd_sc_hd__clkbuf_4 fanout909 (.A(net914),
    .X(net909));
 sky130_fd_sc_hd__clkbuf_4 fanout910 (.A(net912),
    .X(net910));
 sky130_fd_sc_hd__clkbuf_2 fanout911 (.A(net912),
    .X(net911));
 sky130_fd_sc_hd__buf_2 fanout912 (.A(net914),
    .X(net912));
 sky130_fd_sc_hd__buf_4 fanout913 (.A(net914),
    .X(net913));
 sky130_fd_sc_hd__buf_2 fanout914 (.A(net936),
    .X(net914));
 sky130_fd_sc_hd__clkbuf_4 fanout915 (.A(net920),
    .X(net915));
 sky130_fd_sc_hd__clkbuf_4 fanout916 (.A(net920),
    .X(net916));
 sky130_fd_sc_hd__clkbuf_4 fanout917 (.A(net920),
    .X(net917));
 sky130_fd_sc_hd__clkbuf_4 fanout918 (.A(net920),
    .X(net918));
 sky130_fd_sc_hd__clkbuf_2 fanout919 (.A(net920),
    .X(net919));
 sky130_fd_sc_hd__buf_2 fanout920 (.A(net936),
    .X(net920));
 sky130_fd_sc_hd__buf_4 fanout921 (.A(net922),
    .X(net921));
 sky130_fd_sc_hd__clkbuf_4 fanout922 (.A(net924),
    .X(net922));
 sky130_fd_sc_hd__buf_4 fanout923 (.A(net924),
    .X(net923));
 sky130_fd_sc_hd__clkbuf_2 fanout924 (.A(net936),
    .X(net924));
 sky130_fd_sc_hd__clkbuf_4 fanout925 (.A(net929),
    .X(net925));
 sky130_fd_sc_hd__clkbuf_4 fanout926 (.A(net929),
    .X(net926));
 sky130_fd_sc_hd__clkbuf_4 fanout927 (.A(net928),
    .X(net927));
 sky130_fd_sc_hd__clkbuf_4 fanout928 (.A(net929),
    .X(net928));
 sky130_fd_sc_hd__clkbuf_4 fanout929 (.A(net935),
    .X(net929));
 sky130_fd_sc_hd__clkbuf_4 fanout930 (.A(net932),
    .X(net930));
 sky130_fd_sc_hd__clkbuf_4 fanout931 (.A(net932),
    .X(net931));
 sky130_fd_sc_hd__buf_2 fanout932 (.A(net935),
    .X(net932));
 sky130_fd_sc_hd__clkbuf_4 fanout933 (.A(net934),
    .X(net933));
 sky130_fd_sc_hd__clkbuf_4 fanout934 (.A(net935),
    .X(net934));
 sky130_fd_sc_hd__clkbuf_2 fanout935 (.A(net936),
    .X(net935));
 sky130_fd_sc_hd__buf_2 fanout936 (.A(net1043),
    .X(net936));
 sky130_fd_sc_hd__clkbuf_4 fanout937 (.A(net938),
    .X(net937));
 sky130_fd_sc_hd__clkbuf_4 fanout938 (.A(net946),
    .X(net938));
 sky130_fd_sc_hd__clkbuf_4 fanout939 (.A(net941),
    .X(net939));
 sky130_fd_sc_hd__clkbuf_4 fanout940 (.A(net941),
    .X(net940));
 sky130_fd_sc_hd__buf_2 fanout941 (.A(net946),
    .X(net941));
 sky130_fd_sc_hd__clkbuf_4 fanout942 (.A(net946),
    .X(net942));
 sky130_fd_sc_hd__clkbuf_2 fanout943 (.A(net946),
    .X(net943));
 sky130_fd_sc_hd__clkbuf_4 fanout944 (.A(net946),
    .X(net944));
 sky130_fd_sc_hd__clkbuf_2 fanout945 (.A(net946),
    .X(net945));
 sky130_fd_sc_hd__buf_2 fanout946 (.A(net954),
    .X(net946));
 sky130_fd_sc_hd__clkbuf_4 fanout947 (.A(net950),
    .X(net947));
 sky130_fd_sc_hd__clkbuf_4 fanout948 (.A(net950),
    .X(net948));
 sky130_fd_sc_hd__clkbuf_4 fanout949 (.A(net950),
    .X(net949));
 sky130_fd_sc_hd__buf_2 fanout950 (.A(net954),
    .X(net950));
 sky130_fd_sc_hd__clkbuf_4 fanout951 (.A(net952),
    .X(net951));
 sky130_fd_sc_hd__clkbuf_4 fanout952 (.A(net953),
    .X(net952));
 sky130_fd_sc_hd__clkbuf_4 fanout953 (.A(net954),
    .X(net953));
 sky130_fd_sc_hd__buf_2 fanout954 (.A(net1043),
    .X(net954));
 sky130_fd_sc_hd__clkbuf_4 fanout955 (.A(net957),
    .X(net955));
 sky130_fd_sc_hd__buf_2 fanout956 (.A(net957),
    .X(net956));
 sky130_fd_sc_hd__clkbuf_4 fanout957 (.A(net975),
    .X(net957));
 sky130_fd_sc_hd__clkbuf_4 fanout958 (.A(net959),
    .X(net958));
 sky130_fd_sc_hd__clkbuf_4 fanout959 (.A(net975),
    .X(net959));
 sky130_fd_sc_hd__clkbuf_4 fanout960 (.A(net964),
    .X(net960));
 sky130_fd_sc_hd__clkbuf_4 fanout961 (.A(net964),
    .X(net961));
 sky130_fd_sc_hd__clkbuf_4 fanout962 (.A(net964),
    .X(net962));
 sky130_fd_sc_hd__clkbuf_4 fanout963 (.A(net964),
    .X(net963));
 sky130_fd_sc_hd__clkbuf_2 fanout964 (.A(net975),
    .X(net964));
 sky130_fd_sc_hd__clkbuf_4 fanout965 (.A(net967),
    .X(net965));
 sky130_fd_sc_hd__clkbuf_2 fanout966 (.A(net967),
    .X(net966));
 sky130_fd_sc_hd__clkbuf_4 fanout967 (.A(net969),
    .X(net967));
 sky130_fd_sc_hd__clkbuf_4 fanout968 (.A(net969),
    .X(net968));
 sky130_fd_sc_hd__clkbuf_2 fanout969 (.A(net975),
    .X(net969));
 sky130_fd_sc_hd__clkbuf_4 fanout970 (.A(net972),
    .X(net970));
 sky130_fd_sc_hd__clkbuf_4 fanout971 (.A(net972),
    .X(net971));
 sky130_fd_sc_hd__buf_2 fanout972 (.A(net975),
    .X(net972));
 sky130_fd_sc_hd__clkbuf_4 fanout973 (.A(net974),
    .X(net973));
 sky130_fd_sc_hd__clkbuf_2 fanout974 (.A(net975),
    .X(net974));
 sky130_fd_sc_hd__clkbuf_4 fanout975 (.A(net1043),
    .X(net975));
 sky130_fd_sc_hd__clkbuf_4 fanout976 (.A(net977),
    .X(net976));
 sky130_fd_sc_hd__clkbuf_4 fanout977 (.A(net998),
    .X(net977));
 sky130_fd_sc_hd__clkbuf_4 fanout978 (.A(net980),
    .X(net978));
 sky130_fd_sc_hd__clkbuf_4 fanout979 (.A(net980),
    .X(net979));
 sky130_fd_sc_hd__clkbuf_2 fanout980 (.A(net998),
    .X(net980));
 sky130_fd_sc_hd__clkbuf_4 fanout981 (.A(net984),
    .X(net981));
 sky130_fd_sc_hd__buf_2 fanout982 (.A(net984),
    .X(net982));
 sky130_fd_sc_hd__clkbuf_4 fanout983 (.A(net984),
    .X(net983));
 sky130_fd_sc_hd__clkbuf_2 fanout984 (.A(net998),
    .X(net984));
 sky130_fd_sc_hd__clkbuf_4 fanout985 (.A(net987),
    .X(net985));
 sky130_fd_sc_hd__clkbuf_4 fanout986 (.A(net987),
    .X(net986));
 sky130_fd_sc_hd__buf_2 fanout987 (.A(net998),
    .X(net987));
 sky130_fd_sc_hd__clkbuf_4 fanout988 (.A(net989),
    .X(net988));
 sky130_fd_sc_hd__clkbuf_2 fanout989 (.A(net998),
    .X(net989));
 sky130_fd_sc_hd__clkbuf_4 fanout990 (.A(net992),
    .X(net990));
 sky130_fd_sc_hd__clkbuf_2 fanout991 (.A(net992),
    .X(net991));
 sky130_fd_sc_hd__clkbuf_4 fanout992 (.A(net998),
    .X(net992));
 sky130_fd_sc_hd__clkbuf_4 fanout993 (.A(net994),
    .X(net993));
 sky130_fd_sc_hd__buf_2 fanout994 (.A(net998),
    .X(net994));
 sky130_fd_sc_hd__clkbuf_4 fanout995 (.A(net997),
    .X(net995));
 sky130_fd_sc_hd__clkbuf_4 fanout996 (.A(net997),
    .X(net996));
 sky130_fd_sc_hd__clkbuf_4 fanout997 (.A(net998),
    .X(net997));
 sky130_fd_sc_hd__clkbuf_4 fanout998 (.A(net1041),
    .X(net998));
 sky130_fd_sc_hd__clkbuf_4 fanout999 (.A(net1002),
    .X(net999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(net426),
    .X(net1709));
 sky130_fd_sc_hd__dlygate4sd3_1 hold100 (.A(net436),
    .X(net1799));
 sky130_fd_sc_hd__dlygate4sd3_1 hold101 (.A(net1800),
    .X(reg_rdata[26]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold102 (.A(\u_glbl_reg.reg_rdata[23] ),
    .X(net1801));
 sky130_fd_sc_hd__dlygate4sd3_1 hold103 (.A(net433),
    .X(net1802));
 sky130_fd_sc_hd__dlygate4sd3_1 hold104 (.A(net1803),
    .X(reg_rdata[23]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold105 (.A(\u_glbl_reg.reg_rdata[21] ),
    .X(net1804));
 sky130_fd_sc_hd__dlygate4sd3_1 hold106 (.A(net431),
    .X(net1805));
 sky130_fd_sc_hd__dlygate4sd3_1 hold107 (.A(net1806),
    .X(reg_rdata[21]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold108 (.A(\u_ws281x.reg_rdata[27] ),
    .X(net1807));
 sky130_fd_sc_hd__dlygate4sd3_1 hold109 (.A(_03664_),
    .X(net1808));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(net1710),
    .X(reg_rdata[17]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold110 (.A(net437),
    .X(net1809));
 sky130_fd_sc_hd__dlygate4sd3_1 hold111 (.A(net1810),
    .X(reg_rdata[27]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold112 (.A(\u_glbl_reg.reg_rdata[20] ),
    .X(net1811));
 sky130_fd_sc_hd__dlygate4sd3_1 hold113 (.A(net430),
    .X(net1812));
 sky130_fd_sc_hd__dlygate4sd3_1 hold114 (.A(net1813),
    .X(reg_rdata[20]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold115 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[0].u_bit_reg.data_out ),
    .X(net1814));
 sky130_fd_sc_hd__dlygate4sd3_1 hold116 (.A(\u_gpio.u_reg.reg_out[0] ),
    .X(net1815));
 sky130_fd_sc_hd__dlygate4sd3_1 hold117 (.A(\u_pwm.u_pwm_1.cfg_pwm_run ),
    .X(net1816));
 sky130_fd_sc_hd__dlygate4sd3_1 hold118 (.A(\u_pwm.u_glbl_reg.reg_out[9] ),
    .X(net1817));
 sky130_fd_sc_hd__dlygate4sd3_1 hold119 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(net1818));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\u_glbl_reg.reg_rdata[13] ),
    .X(net1711));
 sky130_fd_sc_hd__dlygate4sd3_1 hold120 (.A(\u_gpio.u_reg.reg_out[2] ),
    .X(net1819));
 sky130_fd_sc_hd__dlygate4sd3_1 hold121 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[4].u_bit_reg.data_out ),
    .X(net1820));
 sky130_fd_sc_hd__dlygate4sd3_1 hold122 (.A(\u_gpio.u_reg.reg_out[4] ),
    .X(net1821));
 sky130_fd_sc_hd__dlygate4sd3_1 hold123 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[1].u_bit_reg.data_out ),
    .X(net1822));
 sky130_fd_sc_hd__dlygate4sd3_1 hold124 (.A(\u_pwm.u_glbl_reg.reg_out[1] ),
    .X(net1823));
 sky130_fd_sc_hd__dlygate4sd3_1 hold125 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[0].u_bit_reg.data_out ),
    .X(net1824));
 sky130_fd_sc_hd__dlygate4sd3_1 hold126 (.A(\u_pwm.u_glbl_reg.reg_out[0] ),
    .X(net1825));
 sky130_fd_sc_hd__dlygate4sd3_1 hold127 (.A(\u_pwm.u_pwm_2.cfg_pwm_run ),
    .X(net1826));
 sky130_fd_sc_hd__dlygate4sd3_1 hold128 (.A(\u_glbl_reg.u_random.n1[17] ),
    .X(net1827));
 sky130_fd_sc_hd__dlygate4sd3_1 hold129 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[5].u_bit_reg.data_out ),
    .X(net1828));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(net422),
    .X(net1712));
 sky130_fd_sc_hd__dlygate4sd3_1 hold130 (.A(_01695_),
    .X(net1829));
 sky130_fd_sc_hd__dlygate4sd3_1 hold131 (.A(\u_gpio.u_reg.reg_out[5] ),
    .X(net1830));
 sky130_fd_sc_hd__dlygate4sd3_1 hold132 (.A(\u_gpio.u_bit[3].u_dglitch.gpio_reg ),
    .X(net1831));
 sky130_fd_sc_hd__dlygate4sd3_1 hold133 (.A(_01689_),
    .X(net1832));
 sky130_fd_sc_hd__dlygate4sd3_1 hold134 (.A(\u_gpio.u_reg.reg_out[3] ),
    .X(net1833));
 sky130_fd_sc_hd__dlygate4sd3_1 hold135 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(net1834));
 sky130_fd_sc_hd__dlygate4sd3_1 hold136 (.A(\u_pwm.u_glbl_reg.reg_out[2] ),
    .X(net1835));
 sky130_fd_sc_hd__dlygate4sd3_1 hold137 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[7].u_bit_reg.data_out ),
    .X(net1836));
 sky130_fd_sc_hd__dlygate4sd3_1 hold138 (.A(_01702_),
    .X(net1837));
 sky130_fd_sc_hd__dlygate4sd3_1 hold139 (.A(\u_gpio.u_reg.reg_out[7] ),
    .X(net1838));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(net1713),
    .X(reg_rdata[13]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold140 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[28].u_bit_reg.data_out ),
    .X(net1839));
 sky130_fd_sc_hd__dlygate4sd3_1 hold141 (.A(_01770_),
    .X(net1840));
 sky130_fd_sc_hd__dlygate4sd3_1 hold142 (.A(_01771_),
    .X(net1841));
 sky130_fd_sc_hd__dlygate4sd3_1 hold143 (.A(\u_gpio.u_reg.reg_out[28] ),
    .X(net1842));
 sky130_fd_sc_hd__dlygate4sd3_1 hold144 (.A(\u_prst_sync.in_data_2s ),
    .X(net1843));
 sky130_fd_sc_hd__dlygate4sd3_1 hold145 (.A(\u_gpio.u_bit[1].u_dglitch.gpio_reg ),
    .X(net1844));
 sky130_fd_sc_hd__dlygate4sd3_1 hold146 (.A(_01682_),
    .X(net1845));
 sky130_fd_sc_hd__dlygate4sd3_1 hold147 (.A(\u_gpio.u_reg.reg_out[1] ),
    .X(net1846));
 sky130_fd_sc_hd__dlygate4sd3_1 hold148 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[6].u_bit_reg.data_out ),
    .X(net1847));
 sky130_fd_sc_hd__dlygate4sd3_1 hold149 (.A(_01699_),
    .X(net1848));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\u_glbl_reg.reg_rdata[18] ),
    .X(net1714));
 sky130_fd_sc_hd__dlygate4sd3_1 hold150 (.A(\u_gpio.u_reg.reg_out[6] ),
    .X(net1849));
 sky130_fd_sc_hd__dlygate4sd3_1 hold151 (.A(\u_gpio.u_bit[9].u_dglitch.gpio_reg ),
    .X(net1850));
 sky130_fd_sc_hd__dlygate4sd3_1 hold152 (.A(_01709_),
    .X(net1851));
 sky130_fd_sc_hd__dlygate4sd3_1 hold153 (.A(\u_gpio.u_reg.reg_out[9] ),
    .X(net1852));
 sky130_fd_sc_hd__dlygate4sd3_1 hold154 (.A(\u_glbl_reg.u_random.n0[0] ),
    .X(net1853));
 sky130_fd_sc_hd__dlygate4sd3_1 hold155 (.A(\u_glbl_reg.u_random.n1[28] ),
    .X(net1854));
 sky130_fd_sc_hd__dlygate4sd3_1 hold156 (.A(\u_glbl_reg.u_random.n1[31] ),
    .X(net1855));
 sky130_fd_sc_hd__dlygate4sd3_1 hold157 (.A(\u_glbl_reg.u_random.n1[0] ),
    .X(net1856));
 sky130_fd_sc_hd__dlygate4sd3_1 hold158 (.A(\u_glbl_reg.u_random.n1[2] ),
    .X(net1857));
 sky130_fd_sc_hd__dlygate4sd3_1 hold159 (.A(\u_glbl_reg.u_random.n1[4] ),
    .X(net1858));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(net427),
    .X(net1715));
 sky130_fd_sc_hd__dlygate4sd3_1 hold160 (.A(\u_glbl_reg.u_random.n1[23] ),
    .X(net1859));
 sky130_fd_sc_hd__dlygate4sd3_1 hold161 (.A(\u_glbl_reg.u_random.n1[20] ),
    .X(net1860));
 sky130_fd_sc_hd__dlygate4sd3_1 hold162 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[16].u_bit_reg.data_out ),
    .X(net1861));
 sky130_fd_sc_hd__dlygate4sd3_1 hold163 (.A(\u_gpio.u_reg.reg_out[16] ),
    .X(net1862));
 sky130_fd_sc_hd__dlygate4sd3_1 hold164 (.A(\u_glbl_reg.u_random.n1[21] ),
    .X(net1863));
 sky130_fd_sc_hd__dlygate4sd3_1 hold165 (.A(\u_glbl_reg.u_random.n1[12] ),
    .X(net1864));
 sky130_fd_sc_hd__dlygate4sd3_1 hold166 (.A(\u_glbl_reg.u_random.n1[15] ),
    .X(net1865));
 sky130_fd_sc_hd__dlygate4sd3_1 hold167 (.A(\u_glbl_reg.u_random.n1[30] ),
    .X(net1866));
 sky130_fd_sc_hd__dlygate4sd3_1 hold168 (.A(\u_glbl_reg.u_random.n1[9] ),
    .X(net1867));
 sky130_fd_sc_hd__dlygate4sd3_1 hold169 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[8].u_bit_reg.data_out ),
    .X(net1868));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(net1716),
    .X(reg_rdata[18]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold170 (.A(\u_gpio.u_reg.reg_out[8] ),
    .X(net1869));
 sky130_fd_sc_hd__dlygate4sd3_1 hold171 (.A(\u_glbl_reg.u_random.n1[8] ),
    .X(net1870));
 sky130_fd_sc_hd__dlygate4sd3_1 hold172 (.A(\u_glbl_reg.u_random.n1[3] ),
    .X(net1871));
 sky130_fd_sc_hd__dlygate4sd3_1 hold173 (.A(\u_glbl_reg.u_random.n1[19] ),
    .X(net1872));
 sky130_fd_sc_hd__dlygate4sd3_1 hold174 (.A(\u_glbl_reg.u_random.n1[27] ),
    .X(net1873));
 sky130_fd_sc_hd__dlygate4sd3_1 hold175 (.A(\u_glbl_reg.u_random.n0[15] ),
    .X(net1874));
 sky130_fd_sc_hd__dlygate4sd3_1 hold176 (.A(\u_rst_sync.in_data_2s ),
    .X(net1875));
 sky130_fd_sc_hd__dlygate4sd3_1 hold177 (.A(\u_glbl_reg.u_random.n1[24] ),
    .X(net1876));
 sky130_fd_sc_hd__dlygate4sd3_1 hold178 (.A(\u_glbl_reg.u_random.n1[5] ),
    .X(net1877));
 sky130_fd_sc_hd__dlygate4sd3_1 hold179 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[11].u_bit_reg.data_out ),
    .X(net1878));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\u_glbl_reg.reg_rdata[12] ),
    .X(net1717));
 sky130_fd_sc_hd__dlygate4sd3_1 hold180 (.A(\u_gpio.u_reg.reg_out[11] ),
    .X(net1879));
 sky130_fd_sc_hd__dlygate4sd3_1 hold181 (.A(\u_glbl_reg.u_random.n1[11] ),
    .X(net1880));
 sky130_fd_sc_hd__dlygate4sd3_1 hold182 (.A(\u_glbl_reg.u_random.n0[9] ),
    .X(net1881));
 sky130_fd_sc_hd__dlygate4sd3_1 hold183 (.A(\u_glbl_reg.u_random.n1[18] ),
    .X(net1882));
 sky130_fd_sc_hd__dlygate4sd3_1 hold184 (.A(\u_glbl_reg.u_random.n0[2] ),
    .X(net1883));
 sky130_fd_sc_hd__dlygate4sd3_1 hold185 (.A(\u_glbl_reg.u_random.n0[17] ),
    .X(net1884));
 sky130_fd_sc_hd__dlygate4sd3_1 hold186 (.A(\u_glbl_reg.u_random.n1[10] ),
    .X(net1885));
 sky130_fd_sc_hd__dlygate4sd3_1 hold187 (.A(\u_glbl_reg.u_random.n1[29] ),
    .X(net1886));
 sky130_fd_sc_hd__dlygate4sd3_1 hold188 (.A(\u_glbl_reg.u_random.n1[16] ),
    .X(net1887));
 sky130_fd_sc_hd__dlygate4sd3_1 hold189 (.A(\u_glbl_reg.u_random.n1[26] ),
    .X(net1888));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(net421),
    .X(net1718));
 sky130_fd_sc_hd__dlygate4sd3_1 hold190 (.A(\u_glbl_reg.u_random.n0[8] ),
    .X(net1889));
 sky130_fd_sc_hd__dlygate4sd3_1 hold191 (.A(\u_glbl_reg.u_random.n1[14] ),
    .X(net1890));
 sky130_fd_sc_hd__dlygate4sd3_1 hold192 (.A(\u_glbl_reg.u_random.n1[25] ),
    .X(net1891));
 sky130_fd_sc_hd__dlygate4sd3_1 hold193 (.A(\u_glbl_reg.u_random.n0[24] ),
    .X(net1892));
 sky130_fd_sc_hd__dlygate4sd3_1 hold194 (.A(\u_glbl_reg.u_random.n1[22] ),
    .X(net1893));
 sky130_fd_sc_hd__dlygate4sd3_1 hold195 (.A(\u_glbl_reg.u_random.n0[27] ),
    .X(net1894));
 sky130_fd_sc_hd__dlygate4sd3_1 hold196 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[13].u_bit_reg.data_out ),
    .X(net1895));
 sky130_fd_sc_hd__dlygate4sd3_1 hold197 (.A(\u_gpio.u_reg.reg_out[13] ),
    .X(net1896));
 sky130_fd_sc_hd__dlygate4sd3_1 hold198 (.A(\u_glbl_reg.u_random.n0[28] ),
    .X(net1897));
 sky130_fd_sc_hd__dlygate4sd3_1 hold199 (.A(\u_glbl_reg.u_random.n1[13] ),
    .X(net1898));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(net1719),
    .X(reg_rdata[12]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold200 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[12].u_bit_reg.data_out ),
    .X(net1899));
 sky130_fd_sc_hd__dlygate4sd3_1 hold201 (.A(\u_gpio.u_reg.reg_out[12] ),
    .X(net1900));
 sky130_fd_sc_hd__dlygate4sd3_1 hold202 (.A(\u_glbl_reg.u_random.n0[20] ),
    .X(net1901));
 sky130_fd_sc_hd__dlygate4sd3_1 hold203 (.A(\u_glbl_reg.u_random.n1[1] ),
    .X(net1902));
 sky130_fd_sc_hd__dlygate4sd3_1 hold204 (.A(\u_glbl_reg.u_random.n0[30] ),
    .X(net1903));
 sky130_fd_sc_hd__dlygate4sd3_1 hold205 (.A(\u_glbl_reg.u_random.n1[6] ),
    .X(net1904));
 sky130_fd_sc_hd__dlygate4sd3_1 hold206 (.A(\u_glbl_reg.u_random.n0[23] ),
    .X(net1905));
 sky130_fd_sc_hd__dlygate4sd3_1 hold207 (.A(\u_glbl_reg.u_random.n0[4] ),
    .X(net1906));
 sky130_fd_sc_hd__dlygate4sd3_1 hold208 (.A(\u_glbl_reg.u_random.n0[11] ),
    .X(net1907));
 sky130_fd_sc_hd__dlygate4sd3_1 hold209 (.A(\u_glbl_reg.u_random.n0[10] ),
    .X(net1908));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\u_glbl_reg.reg_rdata[15] ),
    .X(net1720));
 sky130_fd_sc_hd__dlygate4sd3_1 hold210 (.A(\u_glbl_reg.u_random.n0[14] ),
    .X(net1909));
 sky130_fd_sc_hd__dlygate4sd3_1 hold211 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[27].u_bit_reg.data_out ),
    .X(net1910));
 sky130_fd_sc_hd__dlygate4sd3_1 hold212 (.A(\u_gpio.u_reg.reg_out[27] ),
    .X(net1911));
 sky130_fd_sc_hd__dlygate4sd3_1 hold213 (.A(\u_glbl_reg.u_random.n0[29] ),
    .X(net1912));
 sky130_fd_sc_hd__dlygate4sd3_1 hold214 (.A(\u_glbl_reg.u_random.n0[31] ),
    .X(net1913));
 sky130_fd_sc_hd__dlygate4sd3_1 hold215 (.A(\u_glbl_reg.u_random.n1[7] ),
    .X(net1914));
 sky130_fd_sc_hd__dlygate4sd3_1 hold216 (.A(\u_glbl_reg.u_random.n0[26] ),
    .X(net1915));
 sky130_fd_sc_hd__dlygate4sd3_1 hold217 (.A(\u_glbl_reg.u_random.n0[3] ),
    .X(net1916));
 sky130_fd_sc_hd__dlygate4sd3_1 hold218 (.A(\u_glbl_reg.u_random.n0[16] ),
    .X(net1917));
 sky130_fd_sc_hd__dlygate4sd3_1 hold219 (.A(\u_glbl_reg.u_random.n0[1] ),
    .X(net1918));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(net424),
    .X(net1721));
 sky130_fd_sc_hd__dlygate4sd3_1 hold220 (.A(\u_glbl_reg.u_random.n0[5] ),
    .X(net1919));
 sky130_fd_sc_hd__dlygate4sd3_1 hold221 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[31].u_bit_reg.data_out ),
    .X(net1920));
 sky130_fd_sc_hd__dlygate4sd3_1 hold222 (.A(\u_gpio.u_reg.reg_out[31] ),
    .X(net1921));
 sky130_fd_sc_hd__dlygate4sd3_1 hold223 (.A(\u_gpio.u_bit[25].u_dglitch.gpio_reg ),
    .X(net1922));
 sky130_fd_sc_hd__dlygate4sd3_1 hold224 (.A(_01760_),
    .X(net1923));
 sky130_fd_sc_hd__dlygate4sd3_1 hold225 (.A(_01761_),
    .X(net1924));
 sky130_fd_sc_hd__dlygate4sd3_1 hold226 (.A(\u_gpio.u_reg.reg_out[25] ),
    .X(net1925));
 sky130_fd_sc_hd__dlygate4sd3_1 hold227 (.A(\u_glbl_reg.u_random.n0[6] ),
    .X(net1926));
 sky130_fd_sc_hd__dlygate4sd3_1 hold228 (.A(\u_glbl_reg.u_random.n0[19] ),
    .X(net1927));
 sky130_fd_sc_hd__dlygate4sd3_1 hold229 (.A(\u_glbl_reg.u_random.n0[22] ),
    .X(net1928));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(net1722),
    .X(reg_rdata[15]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold230 (.A(\u_glbl_reg.u_random.n0[12] ),
    .X(net1929));
 sky130_fd_sc_hd__dlygate4sd3_1 hold231 (.A(\u_glbl_reg.u_random.n0[21] ),
    .X(net1930));
 sky130_fd_sc_hd__dlygate4sd3_1 hold232 (.A(\u_glbl_reg.u_random.n0[18] ),
    .X(net1931));
 sky130_fd_sc_hd__dlygate4sd3_1 hold233 (.A(\u_glbl_reg.u_random.n0[25] ),
    .X(net1932));
 sky130_fd_sc_hd__dlygate4sd3_1 hold234 (.A(\u_gpio.u_bit[14].u_dglitch.gpio_reg ),
    .X(net1933));
 sky130_fd_sc_hd__dlygate4sd3_1 hold235 (.A(_01727_),
    .X(net1934));
 sky130_fd_sc_hd__dlygate4sd3_1 hold236 (.A(_01728_),
    .X(net1935));
 sky130_fd_sc_hd__dlygate4sd3_1 hold237 (.A(\u_gpio.u_reg.reg_out[14] ),
    .X(net1936));
 sky130_fd_sc_hd__dlygate4sd3_1 hold238 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[26].u_bit_reg.data_out ),
    .X(net1937));
 sky130_fd_sc_hd__dlygate4sd3_1 hold239 (.A(\u_gpio.u_reg.reg_out[26] ),
    .X(net1938));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\u_glbl_reg.reg_rdata[11] ),
    .X(net1723));
 sky130_fd_sc_hd__dlygate4sd3_1 hold240 (.A(\u_glbl_reg.u_random.n0[7] ),
    .X(net1939));
 sky130_fd_sc_hd__dlygate4sd3_1 hold241 (.A(\u_glbl_reg.u_random.n0[13] ),
    .X(net1940));
 sky130_fd_sc_hd__dlygate4sd3_1 hold242 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[20].u_bit_reg.data_out ),
    .X(net1941));
 sky130_fd_sc_hd__dlygate4sd3_1 hold243 (.A(\u_gpio.u_reg.reg_out[20] ),
    .X(net1942));
 sky130_fd_sc_hd__dlygate4sd3_1 hold244 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[23].u_bit_reg.data_out ),
    .X(net1943));
 sky130_fd_sc_hd__dlygate4sd3_1 hold245 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[29].u_bit_reg.data_out ),
    .X(net1944));
 sky130_fd_sc_hd__dlygate4sd3_1 hold246 (.A(\u_gpio.u_reg.reg_out[29] ),
    .X(net1945));
 sky130_fd_sc_hd__dlygate4sd3_1 hold247 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[19].u_bit_reg.data_out ),
    .X(net1946));
 sky130_fd_sc_hd__dlygate4sd3_1 hold248 (.A(\u_gpio.u_reg.reg_out[19] ),
    .X(net1947));
 sky130_fd_sc_hd__dlygate4sd3_1 hold249 (.A(\u_pwm.u_pwm_0.cfg_pwm_run ),
    .X(net1948));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(net420),
    .X(net1724));
 sky130_fd_sc_hd__dlygate4sd3_1 hold250 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[24].u_bit_reg.data_out ),
    .X(net1949));
 sky130_fd_sc_hd__dlygate4sd3_1 hold251 (.A(\u_gpio.u_reg.reg_out[24] ),
    .X(net1950));
 sky130_fd_sc_hd__dlygate4sd3_1 hold252 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[18].u_bit_reg.data_out ),
    .X(net1951));
 sky130_fd_sc_hd__dlygate4sd3_1 hold253 (.A(\u_gpio.u_reg.reg_out[18] ),
    .X(net1952));
 sky130_fd_sc_hd__dlygate4sd3_1 hold254 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[15].u_bit_reg.data_out ),
    .X(net1953));
 sky130_fd_sc_hd__dlygate4sd3_1 hold255 (.A(\u_gpio.u_reg.reg_out[15] ),
    .X(net1954));
 sky130_fd_sc_hd__dlygate4sd3_1 hold256 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[21].u_bit_reg.data_out ),
    .X(net1955));
 sky130_fd_sc_hd__dlygate4sd3_1 hold257 (.A(\u_gpio.u_reg.reg_out[21] ),
    .X(net1956));
 sky130_fd_sc_hd__dlygate4sd3_1 hold258 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[17].u_bit_reg.data_out ),
    .X(net1957));
 sky130_fd_sc_hd__dlygate4sd3_1 hold259 (.A(\u_gpio.u_reg.reg_out[17] ),
    .X(net1958));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(net1725),
    .X(reg_rdata[11]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold260 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[8].u_bit_reg.data_out ),
    .X(net1959));
 sky130_fd_sc_hd__dlygate4sd3_1 hold261 (.A(_01941_),
    .X(net1960));
 sky130_fd_sc_hd__dlygate4sd3_1 hold262 (.A(\u_glbl_reg.reg_out[8] ),
    .X(net1961));
 sky130_fd_sc_hd__dlygate4sd3_1 hold263 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[22].u_bit_reg.data_out ),
    .X(net1962));
 sky130_fd_sc_hd__dlygate4sd3_1 hold264 (.A(\u_gpio.u_reg.reg_out[22] ),
    .X(net1963));
 sky130_fd_sc_hd__dlygate4sd3_1 hold265 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[19] ),
    .X(net1964));
 sky130_fd_sc_hd__dlygate4sd3_1 hold266 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[13].u_bit_reg.data_out ),
    .X(net1965));
 sky130_fd_sc_hd__dlygate4sd3_1 hold267 (.A(\u_glbl_reg.reg_out[13] ),
    .X(net1966));
 sky130_fd_sc_hd__dlygate4sd3_1 hold268 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[15].u_bit_reg.data_out ),
    .X(net1967));
 sky130_fd_sc_hd__dlygate4sd3_1 hold269 (.A(_02064_),
    .X(net1968));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\u_glbl_reg.reg_rdata[16] ),
    .X(net1726));
 sky130_fd_sc_hd__dlygate4sd3_1 hold270 (.A(\u_glbl_reg.reg_out[15] ),
    .X(net1969));
 sky130_fd_sc_hd__dlygate4sd3_1 hold271 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[5].u_bit_reg.data_out ),
    .X(net1970));
 sky130_fd_sc_hd__dlygate4sd3_1 hold272 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[20] ),
    .X(net1971));
 sky130_fd_sc_hd__dlygate4sd3_1 hold273 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[22] ),
    .X(net1972));
 sky130_fd_sc_hd__dlygate4sd3_1 hold274 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[21] ),
    .X(net1973));
 sky130_fd_sc_hd__dlygate4sd3_1 hold275 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[16] ),
    .X(net1974));
 sky130_fd_sc_hd__dlygate4sd3_1 hold276 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[18] ),
    .X(net1975));
 sky130_fd_sc_hd__dlygate4sd3_1 hold277 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[3].u_bit_reg.data_out ),
    .X(net1976));
 sky130_fd_sc_hd__dlygate4sd3_1 hold278 (.A(\u_pwm.u_glbl_reg.u_reg_2.gen_bit_reg[4].u_bit_reg.data_out ),
    .X(net1977));
 sky130_fd_sc_hd__dlygate4sd3_1 hold279 (.A(\u_gpio.u_bit[30].u_dglitch.gpio_reg ),
    .X(net1978));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(net425),
    .X(net1727));
 sky130_fd_sc_hd__dlygate4sd3_1 hold280 (.A(_01777_),
    .X(net1979));
 sky130_fd_sc_hd__dlygate4sd3_1 hold281 (.A(_01778_),
    .X(net1980));
 sky130_fd_sc_hd__dlygate4sd3_1 hold282 (.A(\u_gpio.u_reg.reg_out[30] ),
    .X(net1981));
 sky130_fd_sc_hd__dlygate4sd3_1 hold283 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[11].u_bit_reg.data_out ),
    .X(net1982));
 sky130_fd_sc_hd__dlygate4sd3_1 hold284 (.A(\u_glbl_reg.reg_out[11] ),
    .X(net1983));
 sky130_fd_sc_hd__dlygate4sd3_1 hold285 (.A(\u_glbl_reg.u_random.n1_plus_n0[1] ),
    .X(net1984));
 sky130_fd_sc_hd__dlygate4sd3_1 hold286 (.A(_02130_),
    .X(net1985));
 sky130_fd_sc_hd__dlygate4sd3_1 hold287 (.A(\u_glbl_reg.reg_out[19] ),
    .X(net1986));
 sky130_fd_sc_hd__dlygate4sd3_1 hold288 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[23] ),
    .X(net1987));
 sky130_fd_sc_hd__dlygate4sd3_1 hold289 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[4].u_bit_reg.data_out ),
    .X(net1988));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(net1728),
    .X(reg_rdata[16]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold290 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[17] ),
    .X(net1989));
 sky130_fd_sc_hd__dlygate4sd3_1 hold291 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[12].u_bit_reg.data_out ),
    .X(net1990));
 sky130_fd_sc_hd__dlygate4sd3_1 hold292 (.A(_02016_),
    .X(net1991));
 sky130_fd_sc_hd__dlygate4sd3_1 hold293 (.A(\u_glbl_reg.reg_out[12] ),
    .X(net1992));
 sky130_fd_sc_hd__dlygate4sd3_1 hold294 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[14].u_bit_reg.data_out ),
    .X(net1993));
 sky130_fd_sc_hd__dlygate4sd3_1 hold295 (.A(\u_glbl_reg.reg_out[14] ),
    .X(net1994));
 sky130_fd_sc_hd__dlygate4sd3_1 hold296 (.A(\u_glbl_reg.u_random.n1_plus_n0[5] ),
    .X(net1995));
 sky130_fd_sc_hd__dlygate4sd3_1 hold297 (.A(_02203_),
    .X(net1996));
 sky130_fd_sc_hd__dlygate4sd3_1 hold298 (.A(\u_glbl_reg.reg_out[23] ),
    .X(net1997));
 sky130_fd_sc_hd__dlygate4sd3_1 hold299 (.A(\u_gpio.u_bit[10].u_dglitch.gpio_reg ),
    .X(net1998));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\u_glbl_reg.reg_ack ),
    .X(net1702));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\u_pwm.blk_sel[1] ),
    .X(net1729));
 sky130_fd_sc_hd__dlygate4sd3_1 hold300 (.A(_01714_),
    .X(net1999));
 sky130_fd_sc_hd__dlygate4sd3_1 hold301 (.A(\u_gpio.u_reg.reg_out[10] ),
    .X(net2000));
 sky130_fd_sc_hd__dlygate4sd3_1 hold302 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[29].u_bit_reg.data_out ),
    .X(net2001));
 sky130_fd_sc_hd__dlygate4sd3_1 hold303 (.A(\u_glbl_reg.reg_out[29] ),
    .X(net2002));
 sky130_fd_sc_hd__dlygate4sd3_1 hold304 (.A(\u_glbl_reg.u_random.n1_plus_n0[9] ),
    .X(net2003));
 sky130_fd_sc_hd__dlygate4sd3_1 hold305 (.A(_02259_),
    .X(net2004));
 sky130_fd_sc_hd__dlygate4sd3_1 hold306 (.A(\u_glbl_reg.reg_out[26] ),
    .X(net2005));
 sky130_fd_sc_hd__dlygate4sd3_1 hold307 (.A(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[3].u_bit_reg.data_out ),
    .X(net2006));
 sky130_fd_sc_hd__dlygate4sd3_1 hold308 (.A(\u_pwm.u_pwm_1.cfg_pwm_dupdate ),
    .X(net2007));
 sky130_fd_sc_hd__dlygate4sd3_1 hold309 (.A(\u_glbl_reg.u_random.n1_plus_n0[0] ),
    .X(net2008));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(_03531_),
    .X(net1730));
 sky130_fd_sc_hd__dlygate4sd3_1 hold310 (.A(_02111_),
    .X(net2009));
 sky130_fd_sc_hd__dlygate4sd3_1 hold311 (.A(\u_glbl_reg.reg_out[18] ),
    .X(net2010));
 sky130_fd_sc_hd__dlygate4sd3_1 hold312 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[3].u_bit_reg.data_out ),
    .X(net2011));
 sky130_fd_sc_hd__dlygate4sd3_1 hold313 (.A(_01852_),
    .X(net2012));
 sky130_fd_sc_hd__dlygate4sd3_1 hold314 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[5].u_bit_reg.data_out ),
    .X(net2013));
 sky130_fd_sc_hd__dlygate4sd3_1 hold315 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[24].u_bit_reg.data_out ),
    .X(net2014));
 sky130_fd_sc_hd__dlygate4sd3_1 hold316 (.A(\u_glbl_reg.reg_out[24] ),
    .X(net2015));
 sky130_fd_sc_hd__dlygate4sd3_1 hold317 (.A(\u_pwm.u_pwm_0.cfg_pwm_dupdate ),
    .X(net2016));
 sky130_fd_sc_hd__dlygate4sd3_1 hold318 (.A(\u_timer.cfg_timer1[14] ),
    .X(net2017));
 sky130_fd_sc_hd__dlygate4sd3_1 hold319 (.A(\u_glbl_reg.u_random.n1_plus_n0[11] ),
    .X(net2018));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(_03532_),
    .X(net1731));
 sky130_fd_sc_hd__dlygate4sd3_1 hold320 (.A(_02292_),
    .X(net2019));
 sky130_fd_sc_hd__dlygate4sd3_1 hold321 (.A(\u_glbl_reg.reg_out[28] ),
    .X(net2020));
 sky130_fd_sc_hd__dlygate4sd3_1 hold322 (.A(\u_timer.cfg_timer1[9] ),
    .X(net2021));
 sky130_fd_sc_hd__dlygate4sd3_1 hold323 (.A(\u_timer.cfg_timer1[8] ),
    .X(net2022));
 sky130_fd_sc_hd__dlygate4sd3_1 hold324 (.A(\u_timer.cfg_timer1[10] ),
    .X(net2023));
 sky130_fd_sc_hd__dlygate4sd3_1 hold325 (.A(\u_timer.cfg_timer1[11] ),
    .X(net2024));
 sky130_fd_sc_hd__dlygate4sd3_1 hold326 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[22].u_bit_reg.data_out ),
    .X(net2025));
 sky130_fd_sc_hd__dlygate4sd3_1 hold327 (.A(\u_glbl_reg.reg_out[22] ),
    .X(net2026));
 sky130_fd_sc_hd__dlygate4sd3_1 hold328 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[19] ),
    .X(net2027));
 sky130_fd_sc_hd__dlygate4sd3_1 hold329 (.A(\u_glbl_reg.u_random.n1_plus_n0[31] ),
    .X(net2028));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(_03534_),
    .X(net1732));
 sky130_fd_sc_hd__dlygate4sd3_1 hold330 (.A(_02076_),
    .X(net2029));
 sky130_fd_sc_hd__dlygate4sd3_1 hold331 (.A(_02096_),
    .X(net2030));
 sky130_fd_sc_hd__dlygate4sd3_1 hold332 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[9].u_bit_reg.data_out ),
    .X(net2031));
 sky130_fd_sc_hd__dlygate4sd3_1 hold333 (.A(_01958_),
    .X(net2032));
 sky130_fd_sc_hd__dlygate4sd3_1 hold334 (.A(\u_glbl_reg.reg_out[9] ),
    .X(net2033));
 sky130_fd_sc_hd__dlygate4sd3_1 hold335 (.A(\u_timer.cfg_timer1[13] ),
    .X(net2034));
 sky130_fd_sc_hd__dlygate4sd3_1 hold336 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[30].u_bit_reg.data_out ),
    .X(net2035));
 sky130_fd_sc_hd__dlygate4sd3_1 hold337 (.A(\u_glbl_reg.u_random.n1_plus_n0[10] ),
    .X(net2036));
 sky130_fd_sc_hd__dlygate4sd3_1 hold338 (.A(\u_glbl_reg.reg_out[27] ),
    .X(net2037));
 sky130_fd_sc_hd__dlygate4sd3_1 hold339 (.A(\u_timer.cfg_timer1[15] ),
    .X(net2038));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(net447),
    .X(net1733));
 sky130_fd_sc_hd__dlygate4sd3_1 hold340 (.A(\u_timer.cfg_timer1[12] ),
    .X(net2039));
 sky130_fd_sc_hd__dlygate4sd3_1 hold341 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[31] ),
    .X(net2040));
 sky130_fd_sc_hd__dlygate4sd3_1 hold342 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[24] ),
    .X(net2041));
 sky130_fd_sc_hd__dlygate4sd3_1 hold343 (.A(\u_timer.cfg_timer0[7] ),
    .X(net2042));
 sky130_fd_sc_hd__dlygate4sd3_1 hold344 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[26] ),
    .X(net2043));
 sky130_fd_sc_hd__dlygate4sd3_1 hold345 (.A(\u_timer.cfg_timer0[6] ),
    .X(net2044));
 sky130_fd_sc_hd__dlygate4sd3_1 hold346 (.A(\u_timer.cfg_timer0[0] ),
    .X(net2045));
 sky130_fd_sc_hd__dlygate4sd3_1 hold347 (.A(\u_pwm.u_pwm_2.cfg_pwm_dupdate ),
    .X(net2046));
 sky130_fd_sc_hd__dlygate4sd3_1 hold348 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[30] ),
    .X(net2047));
 sky130_fd_sc_hd__dlygate4sd3_1 hold349 (.A(\u_timer.cfg_timer0[4] ),
    .X(net2048));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(net1734),
    .X(reg_rdata[7]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold350 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[25] ),
    .X(net2049));
 sky130_fd_sc_hd__dlygate4sd3_1 hold351 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[10].u_bit_reg.data_out ),
    .X(net2050));
 sky130_fd_sc_hd__dlygate4sd3_1 hold352 (.A(_01979_),
    .X(net2051));
 sky130_fd_sc_hd__dlygate4sd3_1 hold353 (.A(\u_glbl_reg.reg_out[10] ),
    .X(net2052));
 sky130_fd_sc_hd__dlygate4sd3_1 hold354 (.A(\u_timer.cfg_timer0[3] ),
    .X(net2053));
 sky130_fd_sc_hd__dlygate4sd3_1 hold355 (.A(\u_rst_sync.in_data_s ),
    .X(net2054));
 sky130_fd_sc_hd__dlygate4sd3_1 hold356 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[27] ),
    .X(net2055));
 sky130_fd_sc_hd__dlygate4sd3_1 hold357 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[21].u_bit_reg.data_out ),
    .X(net2056));
 sky130_fd_sc_hd__dlygate4sd3_1 hold358 (.A(\u_glbl_reg.reg_out[21] ),
    .X(net2057));
 sky130_fd_sc_hd__dlygate4sd3_1 hold359 (.A(\u_timer.cfg_timer0[5] ),
    .X(net2058));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\u_glbl_reg.reg_rdata[6] ),
    .X(net1735));
 sky130_fd_sc_hd__dlygate4sd3_1 hold360 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[29] ),
    .X(net2059));
 sky130_fd_sc_hd__dlygate4sd3_1 hold361 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[28] ),
    .X(net2060));
 sky130_fd_sc_hd__dlygate4sd3_1 hold362 (.A(\u_timer.cfg_timer0[2] ),
    .X(net2061));
 sky130_fd_sc_hd__dlygate4sd3_1 hold363 (.A(\u_glbl_reg.reg_16[1] ),
    .X(net2062));
 sky130_fd_sc_hd__dlygate4sd3_1 hold364 (.A(\u_glbl_reg.reg_out[1] ),
    .X(net2063));
 sky130_fd_sc_hd__dlygate4sd3_1 hold365 (.A(\u_timer.cfg_timer0[1] ),
    .X(net2064));
 sky130_fd_sc_hd__dlygate4sd3_1 hold366 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[31].u_bit_reg.data_out ),
    .X(net2065));
 sky130_fd_sc_hd__dlygate4sd3_1 hold367 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[16].u_bit_reg.data_out ),
    .X(net2066));
 sky130_fd_sc_hd__dlygate4sd3_1 hold368 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[8] ),
    .X(net2067));
 sky130_fd_sc_hd__dlygate4sd3_1 hold369 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[16] ),
    .X(net2068));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(net446),
    .X(net1736));
 sky130_fd_sc_hd__dlygate4sd3_1 hold370 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[11] ),
    .X(net2069));
 sky130_fd_sc_hd__dlygate4sd3_1 hold371 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[15] ),
    .X(net2070));
 sky130_fd_sc_hd__dlygate4sd3_1 hold372 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[10] ),
    .X(net2071));
 sky130_fd_sc_hd__dlygate4sd3_1 hold373 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[2] ),
    .X(net2072));
 sky130_fd_sc_hd__dlygate4sd3_1 hold374 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[14] ),
    .X(net2073));
 sky130_fd_sc_hd__dlygate4sd3_1 hold375 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[28] ),
    .X(net2074));
 sky130_fd_sc_hd__dlygate4sd3_1 hold376 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[24] ),
    .X(net2075));
 sky130_fd_sc_hd__dlygate4sd3_1 hold377 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[21] ),
    .X(net2076));
 sky130_fd_sc_hd__dlygate4sd3_1 hold378 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[5] ),
    .X(net2077));
 sky130_fd_sc_hd__dlygate4sd3_1 hold379 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[5] ),
    .X(net2078));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(net1737),
    .X(reg_rdata[6]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold380 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[9] ),
    .X(net2079));
 sky130_fd_sc_hd__dlygate4sd3_1 hold381 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[6] ),
    .X(net2080));
 sky130_fd_sc_hd__dlygate4sd3_1 hold382 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[4] ),
    .X(net2081));
 sky130_fd_sc_hd__dlygate4sd3_1 hold383 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[30] ),
    .X(net2082));
 sky130_fd_sc_hd__dlygate4sd3_1 hold384 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[22] ),
    .X(net2083));
 sky130_fd_sc_hd__dlygate4sd3_1 hold385 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[7] ),
    .X(net2084));
 sky130_fd_sc_hd__dlygate4sd3_1 hold386 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[12] ),
    .X(net2085));
 sky130_fd_sc_hd__dlygate4sd3_1 hold387 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[3] ),
    .X(net2086));
 sky130_fd_sc_hd__dlygate4sd3_1 hold388 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[13] ),
    .X(net2087));
 sky130_fd_sc_hd__dlygate4sd3_1 hold389 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[17] ),
    .X(net2088));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\u_glbl_reg.reg_rdata[14] ),
    .X(net1738));
 sky130_fd_sc_hd__dlygate4sd3_1 hold390 (.A(\u_ws281x.u_txd_1.state ),
    .X(net2089));
 sky130_fd_sc_hd__dlygate4sd3_1 hold391 (.A(_03817_),
    .X(net2090));
 sky130_fd_sc_hd__dlygate4sd3_1 hold392 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[6].u_bit_reg.data_out ),
    .X(net2091));
 sky130_fd_sc_hd__dlygate4sd3_1 hold393 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[19] ),
    .X(net2092));
 sky130_fd_sc_hd__dlygate4sd3_1 hold394 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[5] ),
    .X(net2093));
 sky130_fd_sc_hd__dlygate4sd3_1 hold395 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[23] ),
    .X(net2094));
 sky130_fd_sc_hd__dlygate4sd3_1 hold396 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[7] ),
    .X(net2095));
 sky130_fd_sc_hd__dlygate4sd3_1 hold397 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[20] ),
    .X(net2096));
 sky130_fd_sc_hd__dlygate4sd3_1 hold398 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[7].u_bit_reg.data_out ),
    .X(net2097));
 sky130_fd_sc_hd__dlygate4sd3_1 hold399 (.A(_01922_),
    .X(net2098));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(net2347),
    .X(net1703));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(net423),
    .X(net1739));
 sky130_fd_sc_hd__dlygate4sd3_1 hold400 (.A(\u_ws281x.u_txd_0.state ),
    .X(net2099));
 sky130_fd_sc_hd__dlygate4sd3_1 hold401 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[6] ),
    .X(net2100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold402 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[2] ),
    .X(net2101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold403 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[1] ),
    .X(net2102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold404 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[6] ),
    .X(net2103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold405 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[31] ),
    .X(net2104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold406 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[29] ),
    .X(net2105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold407 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[0] ),
    .X(net2106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold408 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[1] ),
    .X(net2107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold409 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[0] ),
    .X(net2108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(net1740),
    .X(reg_rdata[14]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold410 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[18] ),
    .X(net2109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold411 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[11] ),
    .X(net2110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold412 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[13] ),
    .X(net2111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold413 (.A(\u_ws281x.u_reg.reg_2[31] ),
    .X(net2112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold414 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[27] ),
    .X(net2113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold415 (.A(\u_ws281x.u_reg.reg_2[30] ),
    .X(net2114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold416 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[16] ),
    .X(net2115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold417 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[19] ),
    .X(net2116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold418 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[6] ),
    .X(net2117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold419 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[17] ),
    .X(net2118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\u_glbl_reg.reg_rdata[1] ),
    .X(net1741));
 sky130_fd_sc_hd__dlygate4sd3_1 hold420 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[15] ),
    .X(net2119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold421 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[25] ),
    .X(net2120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold422 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[25] ),
    .X(net2121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold423 (.A(\u_glbl_reg.u_random.n1_plus_n0[3] ),
    .X(net2122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold424 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[3] ),
    .X(net2123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold425 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[16] ),
    .X(net2124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold426 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[0] ),
    .X(net2125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold427 (.A(\u_pwm.u_pwm_0.u_reg.reg_2[18] ),
    .X(net2126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold428 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[26] ),
    .X(net2127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold429 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[1] ),
    .X(net2128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(net429),
    .X(net1742));
 sky130_fd_sc_hd__dlygate4sd3_1 hold430 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[5] ),
    .X(net2129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold431 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[14] ),
    .X(net2130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold432 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[7] ),
    .X(net2131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold433 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[9] ),
    .X(net2132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold434 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[22] ),
    .X(net2133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold435 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[2] ),
    .X(net2134));
 sky130_fd_sc_hd__dlygate4sd3_1 hold436 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[3] ),
    .X(net2135));
 sky130_fd_sc_hd__dlygate4sd3_1 hold437 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[4] ),
    .X(net2136));
 sky130_fd_sc_hd__dlygate4sd3_1 hold438 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[7] ),
    .X(net2137));
 sky130_fd_sc_hd__dlygate4sd3_1 hold439 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[12] ),
    .X(net2138));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(net1743),
    .X(reg_rdata[1]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold440 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[1] ),
    .X(net2139));
 sky130_fd_sc_hd__dlygate4sd3_1 hold441 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[11] ),
    .X(net2140));
 sky130_fd_sc_hd__dlygate4sd3_1 hold442 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[11] ),
    .X(net2141));
 sky130_fd_sc_hd__dlygate4sd3_1 hold443 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[0] ),
    .X(net2142));
 sky130_fd_sc_hd__dlygate4sd3_1 hold444 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[2] ),
    .X(net2143));
 sky130_fd_sc_hd__dlygate4sd3_1 hold445 (.A(\u_ws281x.u_reg.u_reg_0.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(net2144));
 sky130_fd_sc_hd__dlygate4sd3_1 hold446 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[10] ),
    .X(net2145));
 sky130_fd_sc_hd__dlygate4sd3_1 hold447 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[13] ),
    .X(net2146));
 sky130_fd_sc_hd__dlygate4sd3_1 hold448 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[9] ),
    .X(net2147));
 sky130_fd_sc_hd__dlygate4sd3_1 hold449 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[3] ),
    .X(net2148));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\u_glbl_reg.reg_rdata[0] ),
    .X(net1744));
 sky130_fd_sc_hd__dlygate4sd3_1 hold450 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[11] ),
    .X(net2149));
 sky130_fd_sc_hd__dlygate4sd3_1 hold451 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[8] ),
    .X(net2150));
 sky130_fd_sc_hd__dlygate4sd3_1 hold452 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[0] ),
    .X(net2151));
 sky130_fd_sc_hd__dlygate4sd3_1 hold453 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[4] ),
    .X(net2152));
 sky130_fd_sc_hd__dlygate4sd3_1 hold454 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[4] ),
    .X(net2153));
 sky130_fd_sc_hd__dlygate4sd3_1 hold455 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[2] ),
    .X(net2154));
 sky130_fd_sc_hd__dlygate4sd3_1 hold456 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[7] ),
    .X(net2155));
 sky130_fd_sc_hd__dlygate4sd3_1 hold457 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[21] ),
    .X(net2156));
 sky130_fd_sc_hd__dlygate4sd3_1 hold458 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[1] ),
    .X(net2157));
 sky130_fd_sc_hd__dlygate4sd3_1 hold459 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[29] ),
    .X(net2158));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(net418),
    .X(net1745));
 sky130_fd_sc_hd__dlygate4sd3_1 hold460 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[12] ),
    .X(net2159));
 sky130_fd_sc_hd__dlygate4sd3_1 hold461 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[15] ),
    .X(net2160));
 sky130_fd_sc_hd__dlygate4sd3_1 hold462 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[16] ),
    .X(net2161));
 sky130_fd_sc_hd__dlygate4sd3_1 hold463 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[5] ),
    .X(net2162));
 sky130_fd_sc_hd__dlygate4sd3_1 hold464 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[14] ),
    .X(net2163));
 sky130_fd_sc_hd__dlygate4sd3_1 hold465 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[2] ),
    .X(net2164));
 sky130_fd_sc_hd__dlygate4sd3_1 hold466 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[3] ),
    .X(net2165));
 sky130_fd_sc_hd__dlygate4sd3_1 hold467 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[4] ),
    .X(net2166));
 sky130_fd_sc_hd__dlygate4sd3_1 hold468 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[23] ),
    .X(net2167));
 sky130_fd_sc_hd__dlygate4sd3_1 hold469 (.A(\u_pwm.u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(net2168));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(net1746),
    .X(reg_rdata[0]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold470 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[17] ),
    .X(net2169));
 sky130_fd_sc_hd__dlygate4sd3_1 hold471 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[4] ),
    .X(net2170));
 sky130_fd_sc_hd__dlygate4sd3_1 hold472 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[26] ),
    .X(net2171));
 sky130_fd_sc_hd__dlygate4sd3_1 hold473 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[12] ),
    .X(net2172));
 sky130_fd_sc_hd__dlygate4sd3_1 hold474 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[7] ),
    .X(net2173));
 sky130_fd_sc_hd__dlygate4sd3_1 hold475 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[0] ),
    .X(net2174));
 sky130_fd_sc_hd__dlygate4sd3_1 hold476 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[3] ),
    .X(net2175));
 sky130_fd_sc_hd__dlygate4sd3_1 hold477 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[13] ),
    .X(net2176));
 sky130_fd_sc_hd__dlygate4sd3_1 hold478 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[10] ),
    .X(net2177));
 sky130_fd_sc_hd__dlygate4sd3_1 hold479 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[9] ),
    .X(net2178));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\u_glbl_reg.reg_rdata[2] ),
    .X(net1747));
 sky130_fd_sc_hd__dlygate4sd3_1 hold480 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[6] ),
    .X(net2179));
 sky130_fd_sc_hd__dlygate4sd3_1 hold481 (.A(\u_pwm.u_pwm_1.u_reg.reg_2[8] ),
    .X(net2180));
 sky130_fd_sc_hd__dlygate4sd3_1 hold482 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[14] ),
    .X(net2181));
 sky130_fd_sc_hd__dlygate4sd3_1 hold483 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[1] ),
    .X(net2182));
 sky130_fd_sc_hd__dlygate4sd3_1 hold484 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[8] ),
    .X(net2183));
 sky130_fd_sc_hd__dlygate4sd3_1 hold485 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[2] ),
    .X(net2184));
 sky130_fd_sc_hd__dlygate4sd3_1 hold486 (.A(\u_pwm.u_pwm_2.u_reg.reg_1[6] ),
    .X(net2185));
 sky130_fd_sc_hd__dlygate4sd3_1 hold487 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[8] ),
    .X(net2186));
 sky130_fd_sc_hd__dlygate4sd3_1 hold488 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[7] ),
    .X(net2187));
 sky130_fd_sc_hd__dlygate4sd3_1 hold489 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[24] ),
    .X(net2188));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(net440),
    .X(net1748));
 sky130_fd_sc_hd__dlygate4sd3_1 hold490 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[9] ),
    .X(net2189));
 sky130_fd_sc_hd__dlygate4sd3_1 hold491 (.A(\u_pwm.u_pwm_1.u_pwm.pwm_ovflow_l ),
    .X(net2190));
 sky130_fd_sc_hd__dlygate4sd3_1 hold492 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[31] ),
    .X(net2191));
 sky130_fd_sc_hd__dlygate4sd3_1 hold493 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[27] ),
    .X(net2192));
 sky130_fd_sc_hd__dlygate4sd3_1 hold494 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[6] ),
    .X(net2193));
 sky130_fd_sc_hd__dlygate4sd3_1 hold495 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[17] ),
    .X(net2194));
 sky130_fd_sc_hd__dlygate4sd3_1 hold496 (.A(\u_glbl_reg.i2cm_intr_s ),
    .X(net2195));
 sky130_fd_sc_hd__dlygate4sd3_1 hold497 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[2] ),
    .X(net2196));
 sky130_fd_sc_hd__dlygate4sd3_1 hold498 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[0] ),
    .X(net2197));
 sky130_fd_sc_hd__dlygate4sd3_1 hold499 (.A(\u_glbl_reg.usb_intr_s ),
    .X(net2198));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(net1704),
    .X(reg_ack));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(net1749),
    .X(reg_rdata[2]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold500 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[14] ),
    .X(net2199));
 sky130_fd_sc_hd__dlygate4sd3_1 hold501 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[12] ),
    .X(net2200));
 sky130_fd_sc_hd__dlygate4sd3_1 hold502 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[10] ),
    .X(net2201));
 sky130_fd_sc_hd__dlygate4sd3_1 hold503 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[28] ),
    .X(net2202));
 sky130_fd_sc_hd__dlygate4sd3_1 hold504 (.A(\u_pwm.u_pwm_1.u_reg.reg_out[28] ),
    .X(net2203));
 sky130_fd_sc_hd__dlygate4sd3_1 hold505 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[18] ),
    .X(net2204));
 sky130_fd_sc_hd__dlygate4sd3_1 hold506 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[5] ),
    .X(net2205));
 sky130_fd_sc_hd__dlygate4sd3_1 hold507 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[10] ),
    .X(net2206));
 sky130_fd_sc_hd__dlygate4sd3_1 hold508 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[15] ),
    .X(net2207));
 sky130_fd_sc_hd__dlygate4sd3_1 hold509 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[1] ),
    .X(net2208));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\u_glbl_reg.reg_rdata[3] ),
    .X(net1750));
 sky130_fd_sc_hd__dlygate4sd3_1 hold510 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[19] ),
    .X(net2209));
 sky130_fd_sc_hd__dlygate4sd3_1 hold511 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[18] ),
    .X(net2210));
 sky130_fd_sc_hd__dlygate4sd3_1 hold512 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[0] ),
    .X(net2211));
 sky130_fd_sc_hd__dlygate4sd3_1 hold513 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[15] ),
    .X(net2212));
 sky130_fd_sc_hd__dlygate4sd3_1 hold514 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[23] ),
    .X(net2213));
 sky130_fd_sc_hd__dlygate4sd3_1 hold515 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[30] ),
    .X(net2214));
 sky130_fd_sc_hd__dlygate4sd3_1 hold516 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[6] ),
    .X(net2215));
 sky130_fd_sc_hd__dlygate4sd3_1 hold517 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[20] ),
    .X(net2216));
 sky130_fd_sc_hd__dlygate4sd3_1 hold518 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[13] ),
    .X(net2217));
 sky130_fd_sc_hd__dlygate4sd3_1 hold519 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[3] ),
    .X(net2218));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(net443),
    .X(net1751));
 sky130_fd_sc_hd__dlygate4sd3_1 hold520 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[6] ),
    .X(net2219));
 sky130_fd_sc_hd__dlygate4sd3_1 hold521 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[1] ),
    .X(net2220));
 sky130_fd_sc_hd__dlygate4sd3_1 hold522 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[2] ),
    .X(net2221));
 sky130_fd_sc_hd__dlygate4sd3_1 hold523 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[3] ),
    .X(net2222));
 sky130_fd_sc_hd__dlygate4sd3_1 hold524 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[2].u_bit_reg.data_out ),
    .X(net2223));
 sky130_fd_sc_hd__dlygate4sd3_1 hold525 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[5] ),
    .X(net2224));
 sky130_fd_sc_hd__dlygate4sd3_1 hold526 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[7] ),
    .X(net2225));
 sky130_fd_sc_hd__dlygate4sd3_1 hold527 (.A(\u_pwm.u_pwm_1.u_reg.reg_0[20] ),
    .X(net2226));
 sky130_fd_sc_hd__dlygate4sd3_1 hold528 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[4] ),
    .X(net2227));
 sky130_fd_sc_hd__dlygate4sd3_1 hold529 (.A(\u_timer.cfg_timer2[1] ),
    .X(net2228));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(net1752),
    .X(reg_rdata[3]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold530 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[4] ),
    .X(net2229));
 sky130_fd_sc_hd__dlygate4sd3_1 hold531 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[9] ),
    .X(net2230));
 sky130_fd_sc_hd__dlygate4sd3_1 hold532 (.A(\u_timer.u_reg.reg_0[21] ),
    .X(net2231));
 sky130_fd_sc_hd__dlygate4sd3_1 hold533 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[4] ),
    .X(net2232));
 sky130_fd_sc_hd__dlygate4sd3_1 hold534 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[3] ),
    .X(net2233));
 sky130_fd_sc_hd__dlygate4sd3_1 hold535 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[18] ),
    .X(net2234));
 sky130_fd_sc_hd__dlygate4sd3_1 hold536 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[16] ),
    .X(net2235));
 sky130_fd_sc_hd__dlygate4sd3_1 hold537 (.A(\u_gpio.u_bit[1].u_dglitch.gpio_ss[0] ),
    .X(net2236));
 sky130_fd_sc_hd__dlygate4sd3_1 hold538 (.A(\u_gpio.u_bit[31].u_dglitch.gpio_ss[0] ),
    .X(net2237));
 sky130_fd_sc_hd__dlygate4sd3_1 hold539 (.A(\u_gpio.u_bit[3].u_dglitch.gpio_ss[0] ),
    .X(net2238));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\u_glbl_reg.reg_rdata[4] ),
    .X(net1753));
 sky130_fd_sc_hd__dlygate4sd3_1 hold540 (.A(\u_timer.cfg_timer1[7] ),
    .X(net2239));
 sky130_fd_sc_hd__dlygate4sd3_1 hold541 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[11] ),
    .X(net2240));
 sky130_fd_sc_hd__dlygate4sd3_1 hold542 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[7] ),
    .X(net2241));
 sky130_fd_sc_hd__dlygate4sd3_1 hold543 (.A(\u_timer.cfg_timer1[4] ),
    .X(net2242));
 sky130_fd_sc_hd__dlygate4sd3_1 hold544 (.A(\u_gpio.u_bit[25].u_dglitch.gpio_ss[0] ),
    .X(net2243));
 sky130_fd_sc_hd__dlygate4sd3_1 hold545 (.A(\u_timer.cfg_timer1[5] ),
    .X(net2244));
 sky130_fd_sc_hd__dlygate4sd3_1 hold546 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[15] ),
    .X(net2245));
 sky130_fd_sc_hd__dlygate4sd3_1 hold547 (.A(\u_gpio.u_bit[0].u_dglitch.gpio_ss[0] ),
    .X(net2246));
 sky130_fd_sc_hd__dlygate4sd3_1 hold548 (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.empty ),
    .X(net2247));
 sky130_fd_sc_hd__dlygate4sd3_1 hold549 (.A(_00654_),
    .X(net2248));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(net444),
    .X(net1754));
 sky130_fd_sc_hd__dlygate4sd3_1 hold550 (.A(\u_gpio.u_bit[4].u_dglitch.gpio_ss[0] ),
    .X(net2249));
 sky130_fd_sc_hd__dlygate4sd3_1 hold551 (.A(\u_timer.cfg_timer2[0] ),
    .X(net2250));
 sky130_fd_sc_hd__dlygate4sd3_1 hold552 (.A(\u_timer.cfg_timer2[5] ),
    .X(net2251));
 sky130_fd_sc_hd__dlygate4sd3_1 hold553 (.A(\u_gpio.u_bit[20].u_dglitch.gpio_ss[0] ),
    .X(net2252));
 sky130_fd_sc_hd__dlygate4sd3_1 hold554 (.A(\u_timer.cfg_timer1[3] ),
    .X(net2253));
 sky130_fd_sc_hd__dlygate4sd3_1 hold555 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[0] ),
    .X(net2254));
 sky130_fd_sc_hd__dlygate4sd3_1 hold556 (.A(\u_gpio.u_bit[2].u_dglitch.gpio_ss[0] ),
    .X(net2255));
 sky130_fd_sc_hd__dlygate4sd3_1 hold557 (.A(\u_gpio.u_bit[24].u_dglitch.gpio_ss[0] ),
    .X(net2256));
 sky130_fd_sc_hd__dlygate4sd3_1 hold558 (.A(\u_gpio.u_bit[10].u_dglitch.gpio_ss[0] ),
    .X(net2257));
 sky130_fd_sc_hd__dlygate4sd3_1 hold559 (.A(\u_timer.cfg_timer2[2] ),
    .X(net2258));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(net1755),
    .X(reg_rdata[4]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold560 (.A(\u_timer.u_reg.reg_0[23] ),
    .X(net2259));
 sky130_fd_sc_hd__dlygate4sd3_1 hold561 (.A(\u_gpio.u_bit[14].u_dglitch.gpio_ss[0] ),
    .X(net2260));
 sky130_fd_sc_hd__dlygate4sd3_1 hold562 (.A(\u_timer.cfg_timer1[6] ),
    .X(net2261));
 sky130_fd_sc_hd__dlygate4sd3_1 hold563 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[17] ),
    .X(net2262));
 sky130_fd_sc_hd__dlygate4sd3_1 hold564 (.A(\u_timer.cfg_timer2[6] ),
    .X(net2263));
 sky130_fd_sc_hd__dlygate4sd3_1 hold565 (.A(\u_gpio.u_bit[15].u_dglitch.gpio_ss[0] ),
    .X(net2264));
 sky130_fd_sc_hd__dlygate4sd3_1 hold566 (.A(\u_gpio.u_bit[12].u_dglitch.gpio_ss[0] ),
    .X(net2265));
 sky130_fd_sc_hd__dlygate4sd3_1 hold567 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[5] ),
    .X(net2266));
 sky130_fd_sc_hd__dlygate4sd3_1 hold568 (.A(\u_timer.u_reg.reg_0[15] ),
    .X(net2267));
 sky130_fd_sc_hd__dlygate4sd3_1 hold569 (.A(\u_timer.u_reg.reg_0[14] ),
    .X(net2268));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\u_glbl_reg.reg_rdata[5] ),
    .X(net1756));
 sky130_fd_sc_hd__dlygate4sd3_1 hold570 (.A(\u_timer.cfg_timer2[4] ),
    .X(net2269));
 sky130_fd_sc_hd__dlygate4sd3_1 hold571 (.A(\u_timer.cfg_timer2[7] ),
    .X(net2270));
 sky130_fd_sc_hd__dlygate4sd3_1 hold572 (.A(\u_gpio.u_bit[26].u_dglitch.gpio_ss[0] ),
    .X(net2271));
 sky130_fd_sc_hd__dlygate4sd3_1 hold573 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[13] ),
    .X(net2272));
 sky130_fd_sc_hd__dlygate4sd3_1 hold574 (.A(\u_gpio.u_bit[16].u_dglitch.gpio_ss[0] ),
    .X(net2273));
 sky130_fd_sc_hd__dlygate4sd3_1 hold575 (.A(\u_timer.u_reg.reg_0[16] ),
    .X(net2274));
 sky130_fd_sc_hd__dlygate4sd3_1 hold576 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[10] ),
    .X(net2275));
 sky130_fd_sc_hd__dlygate4sd3_1 hold577 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[22] ),
    .X(net2276));
 sky130_fd_sc_hd__dlygate4sd3_1 hold578 (.A(\u_gpio.u_bit[9].u_dglitch.gpio_ss[0] ),
    .X(net2277));
 sky130_fd_sc_hd__dlygate4sd3_1 hold579 (.A(\u_glbl_reg.reg_17[25] ),
    .X(net2278));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(net445),
    .X(net1757));
 sky130_fd_sc_hd__dlygate4sd3_1 hold580 (.A(\u_glbl_reg.reg_out[25] ),
    .X(net2279));
 sky130_fd_sc_hd__dlygate4sd3_1 hold581 (.A(\u_timer.cfg_timer2[13] ),
    .X(net2280));
 sky130_fd_sc_hd__dlygate4sd3_1 hold582 (.A(\u_gpio.u_bit[18].u_dglitch.gpio_ss[0] ),
    .X(net2281));
 sky130_fd_sc_hd__dlygate4sd3_1 hold583 (.A(\u_gpio.u_bit[22].u_dglitch.gpio_ss[0] ),
    .X(net2282));
 sky130_fd_sc_hd__dlygate4sd3_1 hold584 (.A(\u_gpio.u_bit[19].u_dglitch.gpio_ss[0] ),
    .X(net2283));
 sky130_fd_sc_hd__dlygate4sd3_1 hold585 (.A(\u_timer.u_reg.reg_0[20] ),
    .X(net2284));
 sky130_fd_sc_hd__dlygate4sd3_1 hold586 (.A(\u_gpio.u_bit[13].u_dglitch.gpio_ss[0] ),
    .X(net2285));
 sky130_fd_sc_hd__dlygate4sd3_1 hold587 (.A(\u_gpio.u_bit[29].u_dglitch.gpio_ss[0] ),
    .X(net2286));
 sky130_fd_sc_hd__dlygate4sd3_1 hold588 (.A(\u_gpio.u_bit[17].u_dglitch.gpio_ss[0] ),
    .X(net2287));
 sky130_fd_sc_hd__dlygate4sd3_1 hold589 (.A(\u_timer.cfg_timer2[12] ),
    .X(net2288));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(net1758),
    .X(reg_rdata[5]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold590 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[1] ),
    .X(net2289));
 sky130_fd_sc_hd__dlygate4sd3_1 hold591 (.A(\u_timer.cfg_timer2[8] ),
    .X(net2290));
 sky130_fd_sc_hd__dlygate4sd3_1 hold592 (.A(\u_timer.cfg_timer2[9] ),
    .X(net2291));
 sky130_fd_sc_hd__dlygate4sd3_1 hold593 (.A(\u_timer.u_reg.reg_0[11] ),
    .X(net2292));
 sky130_fd_sc_hd__dlygate4sd3_1 hold594 (.A(\u_glbl_reg.u_reg_1.flag ),
    .X(net2293));
 sky130_fd_sc_hd__dlygate4sd3_1 hold595 (.A(\u_timer.u_reg.reg_0[12] ),
    .X(net2294));
 sky130_fd_sc_hd__dlygate4sd3_1 hold596 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[20] ),
    .X(net2295));
 sky130_fd_sc_hd__dlygate4sd3_1 hold597 (.A(\u_timer.u_reg.reg_0[17] ),
    .X(net2296));
 sky130_fd_sc_hd__dlygate4sd3_1 hold598 (.A(\u_gpio.u_bit[21].u_dglitch.gpio_ss[0] ),
    .X(net2297));
 sky130_fd_sc_hd__dlygate4sd3_1 hold599 (.A(\u_timer.cfg_timer2[10] ),
    .X(net2298));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\u_glbl_reg.cfg_rst_ctrl[1] ),
    .X(net1705));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\u_glbl_reg.reg_rdata[9] ),
    .X(net1759));
 sky130_fd_sc_hd__dlygate4sd3_1 hold600 (.A(\u_gpio.u_bit[28].u_dglitch.gpio_ss[0] ),
    .X(net2299));
 sky130_fd_sc_hd__dlygate4sd3_1 hold601 (.A(\u_gpio.u_bit[30].u_dglitch.gpio_ss[0] ),
    .X(net2300));
 sky130_fd_sc_hd__dlygate4sd3_1 hold602 (.A(\u_timer.u_reg.reg_0[22] ),
    .X(net2301));
 sky130_fd_sc_hd__dlygate4sd3_1 hold603 (.A(\u_ws281x.u_reg.gfifo[1].u_fifo.full ),
    .X(net2302));
 sky130_fd_sc_hd__dlygate4sd3_1 hold604 (.A(\u_gpio.u_bit[27].u_dglitch.gpio_ss[0] ),
    .X(net2303));
 sky130_fd_sc_hd__dlygate4sd3_1 hold605 (.A(\u_gpio.u_reg.u_reg_4.gen_bit_reg[9].u_bit_reg.data_out ),
    .X(net2304));
 sky130_fd_sc_hd__dlygate4sd3_1 hold606 (.A(\u_gpio.u_bit[11].u_dglitch.gpio_ss[0] ),
    .X(net2305));
 sky130_fd_sc_hd__dlygate4sd3_1 hold607 (.A(\u_prst_sync.in_data_s ),
    .X(net2306));
 sky130_fd_sc_hd__dlygate4sd3_1 hold608 (.A(\u_timer.cfg_timer2[3] ),
    .X(net2307));
 sky130_fd_sc_hd__dlygate4sd3_1 hold609 (.A(\u_timer.cfg_timer2[11] ),
    .X(net2308));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(net449),
    .X(net1760));
 sky130_fd_sc_hd__dlygate4sd3_1 hold610 (.A(\u_timer.cfg_timer1[1] ),
    .X(net2309));
 sky130_fd_sc_hd__dlygate4sd3_1 hold611 (.A(\u_timer.cfg_timer0[14] ),
    .X(net2310));
 sky130_fd_sc_hd__dlygate4sd3_1 hold612 (.A(\u_timer.cfg_timer2[15] ),
    .X(net2311));
 sky130_fd_sc_hd__dlygate4sd3_1 hold613 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[8] ),
    .X(net2312));
 sky130_fd_sc_hd__dlygate4sd3_1 hold614 (.A(\u_glbl_reg.rtc_intr_s ),
    .X(net2313));
 sky130_fd_sc_hd__dlygate4sd3_1 hold615 (.A(\u_timer.u_reg.reg_0[13] ),
    .X(net2314));
 sky130_fd_sc_hd__dlygate4sd3_1 hold616 (.A(\u_gpio.u_bit[8].u_dglitch.gpio_ss[0] ),
    .X(net2315));
 sky130_fd_sc_hd__dlygate4sd3_1 hold617 (.A(\u_timer.cfg_timer2[14] ),
    .X(net2316));
 sky130_fd_sc_hd__dlygate4sd3_1 hold618 (.A(\u_glbl_reg.u_reg4.gen_bit_reg[0].u_bit_reg.data_out ),
    .X(net2317));
 sky130_fd_sc_hd__dlygate4sd3_1 hold619 (.A(\u_glbl_reg.reg_out[0] ),
    .X(net2318));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(net1761),
    .X(reg_rdata[9]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold620 (.A(\u_ws281x.cfg_reset_period[12] ),
    .X(net2319));
 sky130_fd_sc_hd__dlygate4sd3_1 hold621 (.A(\u_timer.u_reg.reg_0[29] ),
    .X(net2320));
 sky130_fd_sc_hd__dlygate4sd3_1 hold622 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[12] ),
    .X(net2321));
 sky130_fd_sc_hd__dlygate4sd3_1 hold623 (.A(\u_timer.cfg_timer1[2] ),
    .X(net2322));
 sky130_fd_sc_hd__dlygate4sd3_1 hold624 (.A(\u_timer.cfg_timer0[12] ),
    .X(net2323));
 sky130_fd_sc_hd__dlygate4sd3_1 hold625 (.A(\u_timer.cfg_timer0[8] ),
    .X(net2324));
 sky130_fd_sc_hd__dlygate4sd3_1 hold626 (.A(\u_pwm.u_pwm_1.u_reg.reg_1[14] ),
    .X(net2325));
 sky130_fd_sc_hd__dlygate4sd3_1 hold627 (.A(\u_timer.cfg_timer0[11] ),
    .X(net2326));
 sky130_fd_sc_hd__dlygate4sd3_1 hold628 (.A(\u_timer.u_reg.reg_0[18] ),
    .X(net2327));
 sky130_fd_sc_hd__dlygate4sd3_1 hold629 (.A(\u_timer.cfg_timer0[9] ),
    .X(net2328));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\u_glbl_reg.reg_rdata[10] ),
    .X(net1762));
 sky130_fd_sc_hd__dlygate4sd3_1 hold630 (.A(\u_ws281x.port1_enb ),
    .X(net2329));
 sky130_fd_sc_hd__dlygate4sd3_1 hold631 (.A(\u_timer.cfg_timer1[0] ),
    .X(net2330));
 sky130_fd_sc_hd__dlygate4sd3_1 hold632 (.A(\u_timer.u_reg.reg_0[30] ),
    .X(net2331));
 sky130_fd_sc_hd__dlygate4sd3_1 hold633 (.A(\u_timer.cfg_timer0[13] ),
    .X(net2332));
 sky130_fd_sc_hd__dlygate4sd3_1 hold634 (.A(\u_timer.u_reg.reg_0[28] ),
    .X(net2333));
 sky130_fd_sc_hd__dlygate4sd3_1 hold635 (.A(\u_pwm.u_pwm_2.u_reg.reg_2[21] ),
    .X(net2334));
 sky130_fd_sc_hd__dlygate4sd3_1 hold636 (.A(\u_timer.u_reg.reg_0[10] ),
    .X(net2335));
 sky130_fd_sc_hd__dlygate4sd3_1 hold637 (.A(\u_timer.cfg_timer0[10] ),
    .X(net2336));
 sky130_fd_sc_hd__dlygate4sd3_1 hold638 (.A(\u_timer.cfg_timer0[15] ),
    .X(net2337));
 sky130_fd_sc_hd__dlygate4sd3_1 hold639 (.A(\u_timer.u_reg.reg_0[19] ),
    .X(net2338));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(net419),
    .X(net1763));
 sky130_fd_sc_hd__dlygate4sd3_1 hold640 (.A(\u_pwm.u_pwm_2.u_reg.reg_0[19] ),
    .X(net2339));
 sky130_fd_sc_hd__dlygate4sd3_1 hold641 (.A(\u_pwm.u_pwm_0.u_reg.reg_1[23] ),
    .X(net2340));
 sky130_fd_sc_hd__dlygate4sd3_1 hold642 (.A(\u_pwm.u_pwm_2.u_pwm.pwm_ovflow_l ),
    .X(net2341));
 sky130_fd_sc_hd__dlygate4sd3_1 hold643 (.A(\u_ws281x.u_txd_0.state ),
    .X(net2342));
 sky130_fd_sc_hd__dlygate4sd3_1 hold644 (.A(_00603_),
    .X(net2343));
 sky130_fd_sc_hd__dlygate4sd3_1 hold645 (.A(\u_timer.u_reg.reg_0[27] ),
    .X(net2344));
 sky130_fd_sc_hd__dlygate4sd3_1 hold646 (.A(\u_semaphore.reg_ack ),
    .X(net2345));
 sky130_fd_sc_hd__dlygate4sd3_1 hold647 (.A(_03700_),
    .X(net2346));
 sky130_fd_sc_hd__dlygate4sd3_1 hold648 (.A(net368),
    .X(net2347));
 sky130_fd_sc_hd__dlygate4sd3_1 hold649 (.A(\u_ws281x.u_txd_1.state ),
    .X(net2348));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(net1764),
    .X(reg_rdata[10]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold650 (.A(\u_pwm.u_pwm_0.u_reg.reg_0[6] ),
    .X(net2349));
 sky130_fd_sc_hd__dlygate4sd3_1 hold66 (.A(\u_glbl_reg.reg_rdata[31] ),
    .X(net1765));
 sky130_fd_sc_hd__dlygate4sd3_1 hold67 (.A(net442),
    .X(net1766));
 sky130_fd_sc_hd__dlygate4sd3_1 hold68 (.A(net1767),
    .X(reg_rdata[31]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold69 (.A(\u_glbl_reg.reg_rdata[8] ),
    .X(net1768));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net367),
    .X(net1706));
 sky130_fd_sc_hd__dlygate4sd3_1 hold70 (.A(net448),
    .X(net1769));
 sky130_fd_sc_hd__dlygate4sd3_1 hold71 (.A(net1770),
    .X(reg_rdata[8]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold72 (.A(\u_pwm.reg_rdata_pwm1[30] ),
    .X(net1771));
 sky130_fd_sc_hd__dlygate4sd3_1 hold73 (.A(_03684_),
    .X(net1772));
 sky130_fd_sc_hd__dlygate4sd3_1 hold74 (.A(_03687_),
    .X(net1773));
 sky130_fd_sc_hd__dlygate4sd3_1 hold75 (.A(net441),
    .X(net1774));
 sky130_fd_sc_hd__dlygate4sd3_1 hold76 (.A(net1775),
    .X(reg_rdata[30]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold77 (.A(\u_ws281x.reg_rdata[29] ),
    .X(net1776));
 sky130_fd_sc_hd__dlygate4sd3_1 hold78 (.A(_03676_),
    .X(net1777));
 sky130_fd_sc_hd__dlygate4sd3_1 hold79 (.A(net439),
    .X(net1778));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net1707),
    .X(qspim_rst_n));
 sky130_fd_sc_hd__dlygate4sd3_1 hold80 (.A(net1779),
    .X(reg_rdata[29]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold81 (.A(\u_ws281x.reg_rdata[25] ),
    .X(net1780));
 sky130_fd_sc_hd__dlygate4sd3_1 hold82 (.A(_03652_),
    .X(net1781));
 sky130_fd_sc_hd__dlygate4sd3_1 hold83 (.A(net435),
    .X(net1782));
 sky130_fd_sc_hd__dlygate4sd3_1 hold84 (.A(net1783),
    .X(reg_rdata[25]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold85 (.A(\u_ws281x.reg_rdata[22] ),
    .X(net1784));
 sky130_fd_sc_hd__dlygate4sd3_1 hold86 (.A(_03634_),
    .X(net1785));
 sky130_fd_sc_hd__dlygate4sd3_1 hold87 (.A(net432),
    .X(net1786));
 sky130_fd_sc_hd__dlygate4sd3_1 hold88 (.A(net1787),
    .X(reg_rdata[22]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold89 (.A(\u_glbl_reg.reg_rdata[24] ),
    .X(net1788));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\u_glbl_reg.reg_rdata[17] ),
    .X(net1708));
 sky130_fd_sc_hd__dlygate4sd3_1 hold90 (.A(net434),
    .X(net1789));
 sky130_fd_sc_hd__dlygate4sd3_1 hold91 (.A(net1790),
    .X(reg_rdata[24]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold92 (.A(\u_glbl_reg.reg_rdata[28] ),
    .X(net1791));
 sky130_fd_sc_hd__dlygate4sd3_1 hold93 (.A(net438),
    .X(net1792));
 sky130_fd_sc_hd__dlygate4sd3_1 hold94 (.A(net1793),
    .X(reg_rdata[28]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold95 (.A(\u_ws281x.reg_rdata[19] ),
    .X(net1794));
 sky130_fd_sc_hd__dlygate4sd3_1 hold96 (.A(_03616_),
    .X(net1795));
 sky130_fd_sc_hd__dlygate4sd3_1 hold97 (.A(net428),
    .X(net1796));
 sky130_fd_sc_hd__dlygate4sd3_1 hold98 (.A(net1797),
    .X(reg_rdata[19]));
 sky130_fd_sc_hd__dlygate4sd3_1 hold99 (.A(\u_glbl_reg.reg_rdata[26] ),
    .X(net1798));
 sky130_fd_sc_hd__buf_6 input1 (.A(cfg_strap_pad_ctrl),
    .X(net1));
 sky130_fd_sc_hd__buf_6 input10 (.A(digital_io_in[16]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input100 (.A(reg_wdata[11]),
    .X(net100));
 sky130_fd_sc_hd__clkbuf_1 input101 (.A(reg_wdata[12]),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_1 input102 (.A(reg_wdata[13]),
    .X(net102));
 sky130_fd_sc_hd__clkbuf_1 input103 (.A(reg_wdata[14]),
    .X(net103));
 sky130_fd_sc_hd__clkbuf_1 input104 (.A(reg_wdata[15]),
    .X(net104));
 sky130_fd_sc_hd__clkbuf_1 input105 (.A(reg_wdata[16]),
    .X(net105));
 sky130_fd_sc_hd__clkbuf_1 input106 (.A(reg_wdata[17]),
    .X(net106));
 sky130_fd_sc_hd__buf_6 input107 (.A(reg_wdata[18]),
    .X(net107));
 sky130_fd_sc_hd__buf_4 input108 (.A(reg_wdata[19]),
    .X(net108));
 sky130_fd_sc_hd__clkbuf_4 input109 (.A(reg_wdata[1]),
    .X(net109));
 sky130_fd_sc_hd__buf_6 input11 (.A(digital_io_in[17]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input110 (.A(reg_wdata[20]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 input111 (.A(reg_wdata[21]),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_1 input112 (.A(reg_wdata[22]),
    .X(net112));
 sky130_fd_sc_hd__clkbuf_2 input113 (.A(reg_wdata[23]),
    .X(net113));
 sky130_fd_sc_hd__dlymetal6s2s_1 input114 (.A(reg_wdata[24]),
    .X(net114));
 sky130_fd_sc_hd__dlymetal6s2s_1 input115 (.A(reg_wdata[25]),
    .X(net115));
 sky130_fd_sc_hd__dlymetal6s2s_1 input116 (.A(reg_wdata[26]),
    .X(net116));
 sky130_fd_sc_hd__dlymetal6s2s_1 input117 (.A(reg_wdata[27]),
    .X(net117));
 sky130_fd_sc_hd__dlymetal6s2s_1 input118 (.A(reg_wdata[28]),
    .X(net118));
 sky130_fd_sc_hd__dlymetal6s2s_1 input119 (.A(reg_wdata[29]),
    .X(net119));
 sky130_fd_sc_hd__buf_6 input12 (.A(digital_io_in[18]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_2 input120 (.A(reg_wdata[2]),
    .X(net120));
 sky130_fd_sc_hd__dlymetal6s2s_1 input121 (.A(reg_wdata[30]),
    .X(net121));
 sky130_fd_sc_hd__clkbuf_1 input122 (.A(reg_wdata[31]),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_1 input123 (.A(reg_wdata[3]),
    .X(net123));
 sky130_fd_sc_hd__clkbuf_1 input124 (.A(reg_wdata[4]),
    .X(net124));
 sky130_fd_sc_hd__clkbuf_1 input125 (.A(reg_wdata[5]),
    .X(net125));
 sky130_fd_sc_hd__buf_2 input126 (.A(reg_wdata[6]),
    .X(net126));
 sky130_fd_sc_hd__clkbuf_2 input127 (.A(reg_wdata[7]),
    .X(net127));
 sky130_fd_sc_hd__clkbuf_1 input128 (.A(reg_wdata[8]),
    .X(net128));
 sky130_fd_sc_hd__buf_6 input129 (.A(reg_wdata[9]),
    .X(net129));
 sky130_fd_sc_hd__buf_6 input13 (.A(digital_io_in[19]),
    .X(net13));
 sky130_fd_sc_hd__buf_6 input130 (.A(reg_wr),
    .X(net130));
 sky130_fd_sc_hd__clkbuf_2 input131 (.A(riscv_tdo),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_2 input132 (.A(riscv_tdo_en),
    .X(net132));
 sky130_fd_sc_hd__dlymetal6s2s_1 input133 (.A(rtc_intr),
    .X(net133));
 sky130_fd_sc_hd__dlymetal6s2s_1 input134 (.A(s_reset_n),
    .X(net134));
 sky130_fd_sc_hd__clkbuf_1 input135 (.A(sflash_do[0]),
    .X(net135));
 sky130_fd_sc_hd__clkbuf_1 input136 (.A(sflash_do[1]),
    .X(net136));
 sky130_fd_sc_hd__clkbuf_1 input137 (.A(sflash_do[2]),
    .X(net137));
 sky130_fd_sc_hd__clkbuf_1 input138 (.A(sflash_do[3]),
    .X(net138));
 sky130_fd_sc_hd__buf_4 input139 (.A(sflash_oen[0]),
    .X(net139));
 sky130_fd_sc_hd__clkbuf_4 input14 (.A(digital_io_in[1]),
    .X(net14));
 sky130_fd_sc_hd__buf_4 input140 (.A(sflash_oen[1]),
    .X(net140));
 sky130_fd_sc_hd__buf_4 input141 (.A(sflash_oen[2]),
    .X(net141));
 sky130_fd_sc_hd__buf_4 input142 (.A(sflash_oen[3]),
    .X(net142));
 sky130_fd_sc_hd__clkbuf_1 input143 (.A(sflash_sck),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_1 input144 (.A(sflash_ss[0]),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_1 input145 (.A(sflash_ss[1]),
    .X(net145));
 sky130_fd_sc_hd__clkbuf_1 input146 (.A(sflash_ss[2]),
    .X(net146));
 sky130_fd_sc_hd__clkbuf_1 input147 (.A(sflash_ss[3]),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 input148 (.A(sm_a1),
    .X(net148));
 sky130_fd_sc_hd__clkbuf_2 input149 (.A(sm_a2),
    .X(net149));
 sky130_fd_sc_hd__buf_6 input15 (.A(digital_io_in[20]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input150 (.A(sm_b1),
    .X(net150));
 sky130_fd_sc_hd__clkbuf_1 input151 (.A(sm_b2),
    .X(net151));
 sky130_fd_sc_hd__clkbuf_4 input152 (.A(spim_miso),
    .X(net152));
 sky130_fd_sc_hd__clkbuf_4 input153 (.A(spim_sck),
    .X(net153));
 sky130_fd_sc_hd__clkbuf_4 input154 (.A(spim_ssn[0]),
    .X(net154));
 sky130_fd_sc_hd__clkbuf_4 input155 (.A(spim_ssn[1]),
    .X(net155));
 sky130_fd_sc_hd__buf_2 input156 (.A(spim_ssn[2]),
    .X(net156));
 sky130_fd_sc_hd__clkbuf_4 input157 (.A(spim_ssn[3]),
    .X(net157));
 sky130_fd_sc_hd__buf_2 input158 (.A(spis_miso),
    .X(net158));
 sky130_fd_sc_hd__clkbuf_2 input159 (.A(system_strap[0]),
    .X(net159));
 sky130_fd_sc_hd__buf_6 input16 (.A(digital_io_in[21]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input160 (.A(system_strap[10]),
    .X(net160));
 sky130_fd_sc_hd__clkbuf_2 input161 (.A(system_strap[11]),
    .X(net161));
 sky130_fd_sc_hd__buf_2 input162 (.A(system_strap[12]),
    .X(net162));
 sky130_fd_sc_hd__clkbuf_2 input163 (.A(system_strap[13]),
    .X(net163));
 sky130_fd_sc_hd__buf_2 input164 (.A(system_strap[14]),
    .X(net164));
 sky130_fd_sc_hd__clkbuf_2 input165 (.A(system_strap[15]),
    .X(net165));
 sky130_fd_sc_hd__buf_2 input166 (.A(system_strap[16]),
    .X(net166));
 sky130_fd_sc_hd__clkbuf_1 input167 (.A(system_strap[17]),
    .X(net167));
 sky130_fd_sc_hd__clkbuf_2 input168 (.A(system_strap[18]),
    .X(net168));
 sky130_fd_sc_hd__buf_2 input169 (.A(system_strap[19]),
    .X(net169));
 sky130_fd_sc_hd__clkbuf_4 input17 (.A(digital_io_in[22]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input170 (.A(system_strap[1]),
    .X(net170));
 sky130_fd_sc_hd__buf_2 input171 (.A(system_strap[20]),
    .X(net171));
 sky130_fd_sc_hd__buf_2 input172 (.A(system_strap[21]),
    .X(net172));
 sky130_fd_sc_hd__buf_2 input173 (.A(system_strap[22]),
    .X(net173));
 sky130_fd_sc_hd__buf_2 input174 (.A(system_strap[23]),
    .X(net174));
 sky130_fd_sc_hd__clkbuf_1 input175 (.A(system_strap[24]),
    .X(net175));
 sky130_fd_sc_hd__clkbuf_1 input176 (.A(system_strap[25]),
    .X(net176));
 sky130_fd_sc_hd__clkbuf_1 input177 (.A(system_strap[26]),
    .X(net177));
 sky130_fd_sc_hd__dlymetal6s2s_1 input178 (.A(system_strap[27]),
    .X(net178));
 sky130_fd_sc_hd__dlymetal6s2s_1 input179 (.A(system_strap[28]),
    .X(net179));
 sky130_fd_sc_hd__buf_2 input18 (.A(digital_io_in[23]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input180 (.A(system_strap[29]),
    .X(net180));
 sky130_fd_sc_hd__dlymetal6s2s_1 input181 (.A(system_strap[2]),
    .X(net181));
 sky130_fd_sc_hd__dlymetal6s2s_1 input182 (.A(system_strap[30]),
    .X(net182));
 sky130_fd_sc_hd__clkbuf_2 input183 (.A(system_strap[31]),
    .X(net183));
 sky130_fd_sc_hd__dlymetal6s2s_1 input184 (.A(system_strap[3]),
    .X(net184));
 sky130_fd_sc_hd__dlymetal6s2s_1 input185 (.A(system_strap[4]),
    .X(net185));
 sky130_fd_sc_hd__dlymetal6s2s_1 input186 (.A(system_strap[5]),
    .X(net186));
 sky130_fd_sc_hd__dlymetal6s2s_1 input187 (.A(system_strap[6]),
    .X(net187));
 sky130_fd_sc_hd__dlymetal6s2s_1 input188 (.A(system_strap[7]),
    .X(net188));
 sky130_fd_sc_hd__buf_2 input189 (.A(system_strap[8]),
    .X(net189));
 sky130_fd_sc_hd__clkbuf_4 input19 (.A(digital_io_in[24]),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_2 input190 (.A(system_strap[9]),
    .X(net190));
 sky130_fd_sc_hd__clkbuf_2 input191 (.A(uart_txd[0]),
    .X(net191));
 sky130_fd_sc_hd__clkbuf_4 input192 (.A(uart_txd[1]),
    .X(net192));
 sky130_fd_sc_hd__dlymetal6s2s_1 input193 (.A(uartm_txd),
    .X(net193));
 sky130_fd_sc_hd__clkbuf_1 input194 (.A(usb_dn_o),
    .X(net194));
 sky130_fd_sc_hd__clkbuf_4 input195 (.A(usb_dp_o),
    .X(net195));
 sky130_fd_sc_hd__clkbuf_1 input196 (.A(usb_intr),
    .X(net196));
 sky130_fd_sc_hd__clkbuf_1 input197 (.A(usb_oen),
    .X(net197));
 sky130_fd_sc_hd__buf_6 input198 (.A(wbd_clk_int),
    .X(net198));
 sky130_fd_sc_hd__clkbuf_2 input2 (.A(cpu_clk),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input20 (.A(digital_io_in[25]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_4 input21 (.A(digital_io_in[26]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 input22 (.A(digital_io_in[27]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_1 input23 (.A(digital_io_in[29]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 input24 (.A(digital_io_in[2]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_4 input25 (.A(digital_io_in[30]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 input26 (.A(digital_io_in[31]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 input27 (.A(digital_io_in[32]),
    .X(net27));
 sky130_fd_sc_hd__buf_4 input28 (.A(digital_io_in[33]),
    .X(net28));
 sky130_fd_sc_hd__buf_4 input29 (.A(digital_io_in[34]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_1 input3 (.A(digital_io_in[0]),
    .X(net3));
 sky130_fd_sc_hd__buf_6 input30 (.A(digital_io_in[35]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(digital_io_in[36]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 input32 (.A(digital_io_in[3]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_1 input33 (.A(digital_io_in[4]),
    .X(net33));
 sky130_fd_sc_hd__buf_4 input34 (.A(digital_io_in[5]),
    .X(net34));
 sky130_fd_sc_hd__buf_6 input35 (.A(digital_io_in[6]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(digital_io_in[7]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_1 input37 (.A(digital_io_in[8]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(digital_io_in[9]),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 input39 (.A(e_reset_n),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(digital_io_in[10]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_1 input40 (.A(i2cm_clk_o),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_1 input41 (.A(i2cm_clk_oen),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 input42 (.A(i2cm_data_o),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_1 input43 (.A(i2cm_data_oen),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_1 input44 (.A(i2cm_intr),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_1 input45 (.A(int_pll_clock),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_1 input46 (.A(ir_intr),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_1 input47 (.A(ir_tx),
    .X(net47));
 sky130_fd_sc_hd__dlymetal6s2s_1 input48 (.A(p_reset_n),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_1 input49 (.A(reg_addr[0]),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_1 input5 (.A(digital_io_in[11]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input50 (.A(reg_addr[10]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_1 input51 (.A(reg_addr[1]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 input52 (.A(reg_addr[2]),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 input53 (.A(reg_addr[3]),
    .X(net53));
 sky130_fd_sc_hd__clkbuf_1 input54 (.A(reg_addr[4]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 input55 (.A(reg_addr[5]),
    .X(net55));
 sky130_fd_sc_hd__clkbuf_4 input56 (.A(reg_addr[6]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_1 input57 (.A(reg_addr[7]),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 input58 (.A(reg_addr[8]),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 input59 (.A(reg_addr[9]),
    .X(net59));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(digital_io_in[12]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input60 (.A(reg_be[0]),
    .X(net60));
 sky130_fd_sc_hd__buf_6 input61 (.A(reg_be[1]),
    .X(net61));
 sky130_fd_sc_hd__buf_6 input62 (.A(reg_be[2]),
    .X(net62));
 sky130_fd_sc_hd__buf_6 input63 (.A(reg_be[3]),
    .X(net63));
 sky130_fd_sc_hd__clkbuf_1 input64 (.A(reg_cs),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 input65 (.A(reg_peri_ack),
    .X(net65));
 sky130_fd_sc_hd__dlymetal6s2s_1 input66 (.A(reg_peri_rdata[0]),
    .X(net66));
 sky130_fd_sc_hd__clkbuf_1 input67 (.A(reg_peri_rdata[10]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_1 input68 (.A(reg_peri_rdata[11]),
    .X(net68));
 sky130_fd_sc_hd__clkbuf_1 input69 (.A(reg_peri_rdata[12]),
    .X(net69));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(digital_io_in[13]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input70 (.A(reg_peri_rdata[13]),
    .X(net70));
 sky130_fd_sc_hd__clkbuf_1 input71 (.A(reg_peri_rdata[14]),
    .X(net71));
 sky130_fd_sc_hd__clkbuf_1 input72 (.A(reg_peri_rdata[15]),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_1 input73 (.A(reg_peri_rdata[16]),
    .X(net73));
 sky130_fd_sc_hd__dlymetal6s2s_1 input74 (.A(reg_peri_rdata[17]),
    .X(net74));
 sky130_fd_sc_hd__dlymetal6s2s_1 input75 (.A(reg_peri_rdata[18]),
    .X(net75));
 sky130_fd_sc_hd__clkbuf_1 input76 (.A(reg_peri_rdata[19]),
    .X(net76));
 sky130_fd_sc_hd__dlymetal6s2s_1 input77 (.A(reg_peri_rdata[1]),
    .X(net77));
 sky130_fd_sc_hd__dlymetal6s2s_1 input78 (.A(reg_peri_rdata[20]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_1 input79 (.A(reg_peri_rdata[21]),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 input8 (.A(digital_io_in[14]),
    .X(net8));
 sky130_fd_sc_hd__dlymetal6s2s_1 input80 (.A(reg_peri_rdata[22]),
    .X(net80));
 sky130_fd_sc_hd__clkbuf_1 input81 (.A(reg_peri_rdata[23]),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_1 input82 (.A(reg_peri_rdata[24]),
    .X(net82));
 sky130_fd_sc_hd__clkbuf_1 input83 (.A(reg_peri_rdata[25]),
    .X(net83));
 sky130_fd_sc_hd__clkbuf_1 input84 (.A(reg_peri_rdata[26]),
    .X(net84));
 sky130_fd_sc_hd__clkbuf_1 input85 (.A(reg_peri_rdata[27]),
    .X(net85));
 sky130_fd_sc_hd__clkbuf_1 input86 (.A(reg_peri_rdata[28]),
    .X(net86));
 sky130_fd_sc_hd__clkbuf_1 input87 (.A(reg_peri_rdata[29]),
    .X(net87));
 sky130_fd_sc_hd__dlymetal6s2s_1 input88 (.A(reg_peri_rdata[2]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 input89 (.A(reg_peri_rdata[30]),
    .X(net89));
 sky130_fd_sc_hd__buf_6 input9 (.A(digital_io_in[15]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input90 (.A(reg_peri_rdata[31]),
    .X(net90));
 sky130_fd_sc_hd__dlymetal6s2s_1 input91 (.A(reg_peri_rdata[3]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 input92 (.A(reg_peri_rdata[4]),
    .X(net92));
 sky130_fd_sc_hd__dlymetal6s2s_1 input93 (.A(reg_peri_rdata[5]),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_1 input94 (.A(reg_peri_rdata[6]),
    .X(net94));
 sky130_fd_sc_hd__dlymetal6s2s_1 input95 (.A(reg_peri_rdata[7]),
    .X(net95));
 sky130_fd_sc_hd__clkbuf_1 input96 (.A(reg_peri_rdata[8]),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_1 input97 (.A(reg_peri_rdata[9]),
    .X(net97));
 sky130_fd_sc_hd__clkbuf_4 input98 (.A(reg_wdata[0]),
    .X(net98));
 sky130_fd_sc_hd__buf_6 input99 (.A(reg_wdata[10]),
    .X(net99));
 sky130_fd_sc_hd__buf_4 max_length1313 (.A(net1314),
    .X(net1313));
 sky130_fd_sc_hd__buf_4 max_length1322 (.A(net1321),
    .X(net1322));
 sky130_fd_sc_hd__buf_4 max_length1431 (.A(net1432),
    .X(net1431));
 sky130_fd_sc_hd__buf_4 max_length1548 (.A(net1547),
    .X(net1548));
 sky130_fd_sc_hd__buf_6 max_length1558 (.A(net1557),
    .X(net1558));
 sky130_fd_sc_hd__buf_4 max_length1570 (.A(net1569),
    .X(net1570));
 sky130_fd_sc_hd__clkbuf_2 max_length5 (.A(clknet_0_mclk),
    .X(net1695));
 sky130_fd_sc_hd__buf_4 max_length721 (.A(net720),
    .X(net721));
 sky130_fd_sc_hd__buf_2 output199 (.A(net199),
    .X(cfg_dc_trim[0]));
 sky130_fd_sc_hd__buf_2 output200 (.A(net200),
    .X(cfg_dc_trim[10]));
 sky130_fd_sc_hd__buf_2 output201 (.A(net201),
    .X(cfg_dc_trim[11]));
 sky130_fd_sc_hd__buf_2 output202 (.A(net202),
    .X(cfg_dc_trim[12]));
 sky130_fd_sc_hd__buf_2 output203 (.A(net203),
    .X(cfg_dc_trim[13]));
 sky130_fd_sc_hd__buf_2 output204 (.A(net204),
    .X(cfg_dc_trim[14]));
 sky130_fd_sc_hd__buf_2 output205 (.A(net205),
    .X(cfg_dc_trim[15]));
 sky130_fd_sc_hd__buf_2 output206 (.A(net206),
    .X(cfg_dc_trim[16]));
 sky130_fd_sc_hd__buf_2 output207 (.A(net207),
    .X(cfg_dc_trim[17]));
 sky130_fd_sc_hd__buf_2 output208 (.A(net208),
    .X(cfg_dc_trim[18]));
 sky130_fd_sc_hd__buf_2 output209 (.A(net209),
    .X(cfg_dc_trim[19]));
 sky130_fd_sc_hd__buf_2 output210 (.A(net210),
    .X(cfg_dc_trim[1]));
 sky130_fd_sc_hd__buf_2 output211 (.A(net211),
    .X(cfg_dc_trim[20]));
 sky130_fd_sc_hd__buf_2 output212 (.A(net212),
    .X(cfg_dc_trim[21]));
 sky130_fd_sc_hd__buf_2 output213 (.A(net213),
    .X(cfg_dc_trim[22]));
 sky130_fd_sc_hd__buf_2 output214 (.A(net214),
    .X(cfg_dc_trim[23]));
 sky130_fd_sc_hd__buf_2 output215 (.A(net215),
    .X(cfg_dc_trim[24]));
 sky130_fd_sc_hd__buf_2 output216 (.A(net216),
    .X(cfg_dc_trim[25]));
 sky130_fd_sc_hd__buf_2 output217 (.A(net217),
    .X(cfg_dc_trim[2]));
 sky130_fd_sc_hd__buf_2 output218 (.A(net218),
    .X(cfg_dc_trim[3]));
 sky130_fd_sc_hd__buf_2 output219 (.A(net219),
    .X(cfg_dc_trim[4]));
 sky130_fd_sc_hd__buf_2 output220 (.A(net220),
    .X(cfg_dc_trim[5]));
 sky130_fd_sc_hd__buf_2 output221 (.A(net221),
    .X(cfg_dc_trim[6]));
 sky130_fd_sc_hd__buf_2 output222 (.A(net222),
    .X(cfg_dc_trim[7]));
 sky130_fd_sc_hd__buf_2 output223 (.A(net223),
    .X(cfg_dc_trim[8]));
 sky130_fd_sc_hd__buf_2 output224 (.A(net224),
    .X(cfg_dc_trim[9]));
 sky130_fd_sc_hd__buf_2 output225 (.A(net225),
    .X(cfg_dco_mode));
 sky130_fd_sc_hd__buf_2 output226 (.A(net1108),
    .X(cfg_pll_enb));
 sky130_fd_sc_hd__buf_2 output227 (.A(net227),
    .X(cfg_pll_fed_div[0]));
 sky130_fd_sc_hd__buf_2 output228 (.A(net228),
    .X(cfg_pll_fed_div[1]));
 sky130_fd_sc_hd__buf_2 output229 (.A(net229),
    .X(cfg_pll_fed_div[2]));
 sky130_fd_sc_hd__buf_2 output230 (.A(net230),
    .X(cfg_pll_fed_div[3]));
 sky130_fd_sc_hd__buf_2 output231 (.A(net231),
    .X(cfg_pll_fed_div[4]));
 sky130_fd_sc_hd__buf_2 output232 (.A(net232),
    .X(cfg_riscv_ctrl[0]));
 sky130_fd_sc_hd__buf_2 output233 (.A(net233),
    .X(cfg_riscv_ctrl[10]));
 sky130_fd_sc_hd__buf_2 output234 (.A(net234),
    .X(cfg_riscv_ctrl[11]));
 sky130_fd_sc_hd__buf_2 output235 (.A(net235),
    .X(cfg_riscv_ctrl[12]));
 sky130_fd_sc_hd__buf_2 output236 (.A(net236),
    .X(cfg_riscv_ctrl[13]));
 sky130_fd_sc_hd__buf_2 output237 (.A(net237),
    .X(cfg_riscv_ctrl[14]));
 sky130_fd_sc_hd__buf_2 output238 (.A(net238),
    .X(cfg_riscv_ctrl[15]));
 sky130_fd_sc_hd__buf_2 output239 (.A(net239),
    .X(cfg_riscv_ctrl[1]));
 sky130_fd_sc_hd__buf_2 output240 (.A(net240),
    .X(cfg_riscv_ctrl[2]));
 sky130_fd_sc_hd__buf_2 output241 (.A(net241),
    .X(cfg_riscv_ctrl[3]));
 sky130_fd_sc_hd__buf_2 output242 (.A(net242),
    .X(cfg_riscv_ctrl[4]));
 sky130_fd_sc_hd__buf_2 output243 (.A(net243),
    .X(cfg_riscv_ctrl[5]));
 sky130_fd_sc_hd__buf_2 output244 (.A(net244),
    .X(cfg_riscv_ctrl[6]));
 sky130_fd_sc_hd__buf_2 output245 (.A(net245),
    .X(cfg_riscv_ctrl[7]));
 sky130_fd_sc_hd__buf_2 output246 (.A(net246),
    .X(cfg_riscv_ctrl[8]));
 sky130_fd_sc_hd__buf_2 output247 (.A(net247),
    .X(cfg_riscv_ctrl[9]));
 sky130_fd_sc_hd__buf_2 output248 (.A(net248),
    .X(cpu_core_rst_n[0]));
 sky130_fd_sc_hd__buf_2 output249 (.A(net249),
    .X(cpu_core_rst_n[1]));
 sky130_fd_sc_hd__buf_2 output250 (.A(net250),
    .X(cpu_core_rst_n[2]));
 sky130_fd_sc_hd__buf_2 output251 (.A(net251),
    .X(cpu_core_rst_n[3]));
 sky130_fd_sc_hd__buf_2 output252 (.A(net252),
    .X(cpu_intf_rst_n));
 sky130_fd_sc_hd__buf_2 output253 (.A(net253),
    .X(digital_io_oen[0]));
 sky130_fd_sc_hd__buf_2 output254 (.A(net254),
    .X(digital_io_oen[10]));
 sky130_fd_sc_hd__buf_2 output255 (.A(net255),
    .X(digital_io_oen[11]));
 sky130_fd_sc_hd__buf_2 output256 (.A(net256),
    .X(digital_io_oen[12]));
 sky130_fd_sc_hd__buf_2 output257 (.A(net257),
    .X(digital_io_oen[13]));
 sky130_fd_sc_hd__buf_2 output258 (.A(net258),
    .X(digital_io_oen[14]));
 sky130_fd_sc_hd__buf_2 output259 (.A(net581),
    .X(digital_io_oen[15]));
 sky130_fd_sc_hd__buf_2 output260 (.A(net582),
    .X(digital_io_oen[16]));
 sky130_fd_sc_hd__buf_2 output261 (.A(net536),
    .X(digital_io_oen[17]));
 sky130_fd_sc_hd__buf_2 output262 (.A(net537),
    .X(digital_io_oen[18]));
 sky130_fd_sc_hd__buf_2 output263 (.A(net538),
    .X(digital_io_oen[19]));
 sky130_fd_sc_hd__buf_2 output264 (.A(net264),
    .X(digital_io_oen[1]));
 sky130_fd_sc_hd__buf_2 output265 (.A(net583),
    .X(digital_io_oen[20]));
 sky130_fd_sc_hd__buf_2 output266 (.A(net602),
    .X(digital_io_oen[21]));
 sky130_fd_sc_hd__buf_2 output267 (.A(net267),
    .X(digital_io_oen[22]));
 sky130_fd_sc_hd__buf_2 output268 (.A(net268),
    .X(digital_io_oen[23]));
 sky130_fd_sc_hd__buf_2 output269 (.A(net269),
    .X(digital_io_oen[24]));
 sky130_fd_sc_hd__buf_2 output270 (.A(net270),
    .X(digital_io_oen[25]));
 sky130_fd_sc_hd__buf_2 output271 (.A(net271),
    .X(digital_io_oen[26]));
 sky130_fd_sc_hd__buf_2 output272 (.A(net272),
    .X(digital_io_oen[27]));
 sky130_fd_sc_hd__buf_2 output273 (.A(net273),
    .X(digital_io_oen[28]));
 sky130_fd_sc_hd__buf_2 output274 (.A(net274),
    .X(digital_io_oen[29]));
 sky130_fd_sc_hd__buf_2 output275 (.A(net275),
    .X(digital_io_oen[2]));
 sky130_fd_sc_hd__buf_2 output276 (.A(net276),
    .X(digital_io_oen[30]));
 sky130_fd_sc_hd__buf_2 output277 (.A(net277),
    .X(digital_io_oen[31]));
 sky130_fd_sc_hd__buf_2 output278 (.A(net278),
    .X(digital_io_oen[32]));
 sky130_fd_sc_hd__buf_2 output279 (.A(net279),
    .X(digital_io_oen[33]));
 sky130_fd_sc_hd__buf_2 output280 (.A(net280),
    .X(digital_io_oen[34]));
 sky130_fd_sc_hd__buf_2 output281 (.A(net281),
    .X(digital_io_oen[35]));
 sky130_fd_sc_hd__buf_2 output282 (.A(net282),
    .X(digital_io_oen[36]));
 sky130_fd_sc_hd__buf_2 output283 (.A(net283),
    .X(digital_io_oen[37]));
 sky130_fd_sc_hd__buf_2 output284 (.A(net284),
    .X(digital_io_oen[3]));
 sky130_fd_sc_hd__buf_2 output285 (.A(net285),
    .X(digital_io_oen[4]));
 sky130_fd_sc_hd__buf_2 output286 (.A(net286),
    .X(digital_io_oen[5]));
 sky130_fd_sc_hd__buf_2 output287 (.A(net287),
    .X(digital_io_oen[6]));
 sky130_fd_sc_hd__buf_2 output288 (.A(net288),
    .X(digital_io_oen[7]));
 sky130_fd_sc_hd__buf_2 output289 (.A(net289),
    .X(digital_io_oen[8]));
 sky130_fd_sc_hd__buf_2 output290 (.A(net290),
    .X(digital_io_oen[9]));
 sky130_fd_sc_hd__buf_2 output291 (.A(net291),
    .X(digital_io_out[0]));
 sky130_fd_sc_hd__buf_2 output292 (.A(net292),
    .X(digital_io_out[10]));
 sky130_fd_sc_hd__buf_2 output293 (.A(net293),
    .X(digital_io_out[11]));
 sky130_fd_sc_hd__buf_2 output294 (.A(net294),
    .X(digital_io_out[12]));
 sky130_fd_sc_hd__buf_2 output295 (.A(net295),
    .X(digital_io_out[13]));
 sky130_fd_sc_hd__buf_2 output296 (.A(net529),
    .X(digital_io_out[14]));
 sky130_fd_sc_hd__buf_2 output297 (.A(net297),
    .X(digital_io_out[15]));
 sky130_fd_sc_hd__buf_2 output298 (.A(net565),
    .X(digital_io_out[16]));
 sky130_fd_sc_hd__buf_2 output299 (.A(net530),
    .X(digital_io_out[17]));
 sky130_fd_sc_hd__buf_2 output300 (.A(net531),
    .X(digital_io_out[18]));
 sky130_fd_sc_hd__buf_2 output301 (.A(net527),
    .X(digital_io_out[19]));
 sky130_fd_sc_hd__buf_2 output302 (.A(net302),
    .X(digital_io_out[1]));
 sky130_fd_sc_hd__buf_2 output303 (.A(net532),
    .X(digital_io_out[20]));
 sky130_fd_sc_hd__buf_2 output304 (.A(net566),
    .X(digital_io_out[21]));
 sky130_fd_sc_hd__buf_2 output305 (.A(net305),
    .X(digital_io_out[22]));
 sky130_fd_sc_hd__buf_2 output306 (.A(net306),
    .X(digital_io_out[23]));
 sky130_fd_sc_hd__buf_2 output307 (.A(net307),
    .X(digital_io_out[24]));
 sky130_fd_sc_hd__buf_2 output308 (.A(net308),
    .X(digital_io_out[25]));
 sky130_fd_sc_hd__buf_2 output309 (.A(net309),
    .X(digital_io_out[26]));
 sky130_fd_sc_hd__buf_2 output310 (.A(net310),
    .X(digital_io_out[27]));
 sky130_fd_sc_hd__buf_2 output311 (.A(net1199),
    .X(digital_io_out[28]));
 sky130_fd_sc_hd__buf_2 output312 (.A(net1197),
    .X(digital_io_out[29]));
 sky130_fd_sc_hd__buf_2 output313 (.A(net313),
    .X(digital_io_out[2]));
 sky130_fd_sc_hd__buf_2 output314 (.A(net1195),
    .X(digital_io_out[30]));
 sky130_fd_sc_hd__buf_2 output315 (.A(net1193),
    .X(digital_io_out[31]));
 sky130_fd_sc_hd__buf_2 output316 (.A(net1191),
    .X(digital_io_out[32]));
 sky130_fd_sc_hd__buf_2 output317 (.A(net1189),
    .X(digital_io_out[33]));
 sky130_fd_sc_hd__buf_2 output318 (.A(net1187),
    .X(digital_io_out[34]));
 sky130_fd_sc_hd__buf_2 output319 (.A(net1185),
    .X(digital_io_out[35]));
 sky130_fd_sc_hd__buf_2 output320 (.A(net1183),
    .X(digital_io_out[36]));
 sky130_fd_sc_hd__buf_2 output321 (.A(net321),
    .X(digital_io_out[37]));
 sky130_fd_sc_hd__buf_2 output322 (.A(net322),
    .X(digital_io_out[3]));
 sky130_fd_sc_hd__buf_2 output323 (.A(net323),
    .X(digital_io_out[4]));
 sky130_fd_sc_hd__buf_2 output324 (.A(net324),
    .X(digital_io_out[5]));
 sky130_fd_sc_hd__buf_2 output325 (.A(net325),
    .X(digital_io_out[6]));
 sky130_fd_sc_hd__buf_2 output326 (.A(net528),
    .X(digital_io_out[7]));
 sky130_fd_sc_hd__buf_2 output327 (.A(net327),
    .X(digital_io_out[8]));
 sky130_fd_sc_hd__buf_2 output328 (.A(net328),
    .X(digital_io_out[9]));
 sky130_fd_sc_hd__buf_2 output329 (.A(net329),
    .X(i2cm_clk_i));
 sky130_fd_sc_hd__buf_2 output330 (.A(net330),
    .X(i2cm_data_i));
 sky130_fd_sc_hd__buf_2 output331 (.A(net331),
    .X(i2cm_rst_n));
 sky130_fd_sc_hd__buf_2 output332 (.A(net332),
    .X(ir_rx));
 sky130_fd_sc_hd__buf_2 output333 (.A(net333),
    .X(irq_lines[0]));
 sky130_fd_sc_hd__buf_2 output334 (.A(net334),
    .X(irq_lines[10]));
 sky130_fd_sc_hd__buf_2 output335 (.A(net335),
    .X(irq_lines[11]));
 sky130_fd_sc_hd__buf_2 output336 (.A(net336),
    .X(irq_lines[12]));
 sky130_fd_sc_hd__buf_2 output337 (.A(net337),
    .X(irq_lines[13]));
 sky130_fd_sc_hd__buf_2 output338 (.A(net338),
    .X(irq_lines[14]));
 sky130_fd_sc_hd__buf_2 output339 (.A(net339),
    .X(irq_lines[15]));
 sky130_fd_sc_hd__buf_2 output340 (.A(net340),
    .X(irq_lines[16]));
 sky130_fd_sc_hd__buf_2 output341 (.A(net341),
    .X(irq_lines[17]));
 sky130_fd_sc_hd__buf_2 output342 (.A(net342),
    .X(irq_lines[18]));
 sky130_fd_sc_hd__buf_2 output343 (.A(net343),
    .X(irq_lines[19]));
 sky130_fd_sc_hd__buf_2 output344 (.A(net344),
    .X(irq_lines[1]));
 sky130_fd_sc_hd__buf_2 output345 (.A(net345),
    .X(irq_lines[20]));
 sky130_fd_sc_hd__buf_2 output346 (.A(net346),
    .X(irq_lines[21]));
 sky130_fd_sc_hd__buf_2 output347 (.A(net347),
    .X(irq_lines[22]));
 sky130_fd_sc_hd__buf_2 output348 (.A(net348),
    .X(irq_lines[23]));
 sky130_fd_sc_hd__buf_2 output349 (.A(net349),
    .X(irq_lines[24]));
 sky130_fd_sc_hd__buf_2 output350 (.A(net350),
    .X(irq_lines[25]));
 sky130_fd_sc_hd__buf_2 output351 (.A(net351),
    .X(irq_lines[26]));
 sky130_fd_sc_hd__buf_2 output352 (.A(net352),
    .X(irq_lines[27]));
 sky130_fd_sc_hd__buf_2 output353 (.A(net353),
    .X(irq_lines[28]));
 sky130_fd_sc_hd__buf_2 output354 (.A(net354),
    .X(irq_lines[29]));
 sky130_fd_sc_hd__buf_2 output355 (.A(net355),
    .X(irq_lines[2]));
 sky130_fd_sc_hd__buf_2 output356 (.A(net356),
    .X(irq_lines[30]));
 sky130_fd_sc_hd__buf_2 output357 (.A(net357),
    .X(irq_lines[31]));
 sky130_fd_sc_hd__buf_2 output358 (.A(net358),
    .X(irq_lines[3]));
 sky130_fd_sc_hd__buf_2 output359 (.A(net359),
    .X(irq_lines[4]));
 sky130_fd_sc_hd__buf_2 output360 (.A(net360),
    .X(irq_lines[5]));
 sky130_fd_sc_hd__buf_2 output361 (.A(net361),
    .X(irq_lines[6]));
 sky130_fd_sc_hd__buf_2 output362 (.A(net362),
    .X(irq_lines[7]));
 sky130_fd_sc_hd__buf_2 output363 (.A(net363),
    .X(irq_lines[8]));
 sky130_fd_sc_hd__buf_2 output364 (.A(net364),
    .X(irq_lines[9]));
 sky130_fd_sc_hd__buf_2 output365 (.A(net1206),
    .X(pll_ref_clk));
 sky130_fd_sc_hd__buf_2 output366 (.A(net533),
    .X(pulse1m_mclk));
 sky130_fd_sc_hd__buf_2 output367 (.A(net1706),
    .X(net1707));
 sky130_fd_sc_hd__buf_2 output368 (.A(net1703),
    .X(net1704));
 sky130_fd_sc_hd__buf_2 output369 (.A(net369),
    .X(reg_peri_addr[0]));
 sky130_fd_sc_hd__buf_2 output370 (.A(net370),
    .X(reg_peri_addr[10]));
 sky130_fd_sc_hd__buf_2 output371 (.A(net371),
    .X(reg_peri_addr[1]));
 sky130_fd_sc_hd__buf_2 output372 (.A(net372),
    .X(reg_peri_addr[2]));
 sky130_fd_sc_hd__buf_2 output373 (.A(net373),
    .X(reg_peri_addr[3]));
 sky130_fd_sc_hd__buf_2 output374 (.A(net374),
    .X(reg_peri_addr[4]));
 sky130_fd_sc_hd__buf_2 output375 (.A(net375),
    .X(reg_peri_addr[5]));
 sky130_fd_sc_hd__buf_2 output376 (.A(net376),
    .X(reg_peri_addr[6]));
 sky130_fd_sc_hd__buf_2 output377 (.A(net377),
    .X(reg_peri_addr[7]));
 sky130_fd_sc_hd__buf_2 output378 (.A(net378),
    .X(reg_peri_addr[8]));
 sky130_fd_sc_hd__buf_2 output379 (.A(net379),
    .X(reg_peri_addr[9]));
 sky130_fd_sc_hd__buf_2 output380 (.A(net380),
    .X(reg_peri_be[0]));
 sky130_fd_sc_hd__buf_2 output381 (.A(net381),
    .X(reg_peri_be[1]));
 sky130_fd_sc_hd__buf_2 output382 (.A(net382),
    .X(reg_peri_be[2]));
 sky130_fd_sc_hd__buf_2 output383 (.A(net383),
    .X(reg_peri_be[3]));
 sky130_fd_sc_hd__buf_2 output384 (.A(net384),
    .X(reg_peri_cs));
 sky130_fd_sc_hd__buf_2 output385 (.A(net385),
    .X(reg_peri_wdata[0]));
 sky130_fd_sc_hd__buf_2 output386 (.A(net386),
    .X(reg_peri_wdata[10]));
 sky130_fd_sc_hd__buf_2 output387 (.A(net387),
    .X(reg_peri_wdata[11]));
 sky130_fd_sc_hd__buf_2 output388 (.A(net388),
    .X(reg_peri_wdata[12]));
 sky130_fd_sc_hd__buf_2 output389 (.A(net389),
    .X(reg_peri_wdata[13]));
 sky130_fd_sc_hd__buf_2 output390 (.A(net390),
    .X(reg_peri_wdata[14]));
 sky130_fd_sc_hd__buf_2 output391 (.A(net391),
    .X(reg_peri_wdata[15]));
 sky130_fd_sc_hd__buf_2 output392 (.A(net392),
    .X(reg_peri_wdata[16]));
 sky130_fd_sc_hd__buf_2 output393 (.A(net393),
    .X(reg_peri_wdata[17]));
 sky130_fd_sc_hd__buf_2 output394 (.A(net394),
    .X(reg_peri_wdata[18]));
 sky130_fd_sc_hd__buf_2 output395 (.A(net395),
    .X(reg_peri_wdata[19]));
 sky130_fd_sc_hd__buf_2 output396 (.A(net396),
    .X(reg_peri_wdata[1]));
 sky130_fd_sc_hd__buf_2 output397 (.A(net397),
    .X(reg_peri_wdata[20]));
 sky130_fd_sc_hd__buf_2 output398 (.A(net398),
    .X(reg_peri_wdata[21]));
 sky130_fd_sc_hd__buf_2 output399 (.A(net399),
    .X(reg_peri_wdata[22]));
 sky130_fd_sc_hd__buf_2 output400 (.A(net400),
    .X(reg_peri_wdata[23]));
 sky130_fd_sc_hd__buf_2 output401 (.A(net401),
    .X(reg_peri_wdata[24]));
 sky130_fd_sc_hd__buf_2 output402 (.A(net402),
    .X(reg_peri_wdata[25]));
 sky130_fd_sc_hd__buf_2 output403 (.A(net403),
    .X(reg_peri_wdata[26]));
 sky130_fd_sc_hd__buf_2 output404 (.A(net404),
    .X(reg_peri_wdata[27]));
 sky130_fd_sc_hd__buf_2 output405 (.A(net405),
    .X(reg_peri_wdata[28]));
 sky130_fd_sc_hd__buf_2 output406 (.A(net406),
    .X(reg_peri_wdata[29]));
 sky130_fd_sc_hd__buf_2 output407 (.A(net407),
    .X(reg_peri_wdata[2]));
 sky130_fd_sc_hd__buf_2 output408 (.A(net408),
    .X(reg_peri_wdata[30]));
 sky130_fd_sc_hd__buf_2 output409 (.A(net409),
    .X(reg_peri_wdata[31]));
 sky130_fd_sc_hd__buf_2 output410 (.A(net410),
    .X(reg_peri_wdata[3]));
 sky130_fd_sc_hd__buf_2 output411 (.A(net411),
    .X(reg_peri_wdata[4]));
 sky130_fd_sc_hd__buf_2 output412 (.A(net412),
    .X(reg_peri_wdata[5]));
 sky130_fd_sc_hd__buf_2 output413 (.A(net413),
    .X(reg_peri_wdata[6]));
 sky130_fd_sc_hd__buf_2 output414 (.A(net414),
    .X(reg_peri_wdata[7]));
 sky130_fd_sc_hd__buf_2 output415 (.A(net415),
    .X(reg_peri_wdata[8]));
 sky130_fd_sc_hd__buf_2 output416 (.A(net416),
    .X(reg_peri_wdata[9]));
 sky130_fd_sc_hd__buf_2 output417 (.A(net417),
    .X(reg_peri_wr));
 sky130_fd_sc_hd__buf_2 output418 (.A(net1745),
    .X(net1746));
 sky130_fd_sc_hd__buf_2 output419 (.A(net1763),
    .X(net1764));
 sky130_fd_sc_hd__buf_2 output420 (.A(net1724),
    .X(net1725));
 sky130_fd_sc_hd__buf_2 output421 (.A(net1718),
    .X(net1719));
 sky130_fd_sc_hd__buf_2 output422 (.A(net1712),
    .X(net1713));
 sky130_fd_sc_hd__buf_2 output423 (.A(net1739),
    .X(net1740));
 sky130_fd_sc_hd__buf_2 output424 (.A(net1721),
    .X(net1722));
 sky130_fd_sc_hd__buf_2 output425 (.A(net1727),
    .X(net1728));
 sky130_fd_sc_hd__buf_2 output426 (.A(net1709),
    .X(net1710));
 sky130_fd_sc_hd__buf_2 output427 (.A(net1715),
    .X(net1716));
 sky130_fd_sc_hd__buf_2 output428 (.A(net1796),
    .X(net1797));
 sky130_fd_sc_hd__buf_2 output429 (.A(net1742),
    .X(net1743));
 sky130_fd_sc_hd__buf_2 output430 (.A(net1812),
    .X(net1813));
 sky130_fd_sc_hd__buf_2 output431 (.A(net1805),
    .X(net1806));
 sky130_fd_sc_hd__buf_2 output432 (.A(net1786),
    .X(net1787));
 sky130_fd_sc_hd__buf_2 output433 (.A(net1802),
    .X(net1803));
 sky130_fd_sc_hd__buf_2 output434 (.A(net1789),
    .X(net1790));
 sky130_fd_sc_hd__buf_2 output435 (.A(net1782),
    .X(net1783));
 sky130_fd_sc_hd__buf_2 output436 (.A(net1799),
    .X(net1800));
 sky130_fd_sc_hd__buf_2 output437 (.A(net1809),
    .X(net1810));
 sky130_fd_sc_hd__buf_2 output438 (.A(net1792),
    .X(net1793));
 sky130_fd_sc_hd__buf_2 output439 (.A(net1778),
    .X(net1779));
 sky130_fd_sc_hd__buf_2 output440 (.A(net1748),
    .X(net1749));
 sky130_fd_sc_hd__buf_2 output441 (.A(net1774),
    .X(net1775));
 sky130_fd_sc_hd__buf_2 output442 (.A(net1766),
    .X(net1767));
 sky130_fd_sc_hd__buf_2 output443 (.A(net1751),
    .X(net1752));
 sky130_fd_sc_hd__buf_2 output444 (.A(net1754),
    .X(net1755));
 sky130_fd_sc_hd__buf_2 output445 (.A(net1757),
    .X(net1758));
 sky130_fd_sc_hd__buf_2 output446 (.A(net1736),
    .X(net1737));
 sky130_fd_sc_hd__buf_2 output447 (.A(net1733),
    .X(net1734));
 sky130_fd_sc_hd__buf_2 output448 (.A(net1769),
    .X(net1770));
 sky130_fd_sc_hd__buf_2 output449 (.A(net1760),
    .X(net1761));
 sky130_fd_sc_hd__buf_2 output450 (.A(net450),
    .X(riscv_tck));
 sky130_fd_sc_hd__buf_2 output451 (.A(net451),
    .X(riscv_tdi));
 sky130_fd_sc_hd__buf_2 output452 (.A(net452),
    .X(riscv_tms));
 sky130_fd_sc_hd__buf_2 output453 (.A(net453),
    .X(riscv_trst_n));
 sky130_fd_sc_hd__clkbuf_1 output454 (.A(net1697),
    .X(rtc_clk));
 sky130_fd_sc_hd__buf_2 output455 (.A(net455),
    .X(sflash_di[0]));
 sky130_fd_sc_hd__buf_2 output456 (.A(net456),
    .X(sflash_di[1]));
 sky130_fd_sc_hd__buf_2 output457 (.A(net457),
    .X(sflash_di[2]));
 sky130_fd_sc_hd__buf_2 output458 (.A(net458),
    .X(sflash_di[3]));
 sky130_fd_sc_hd__buf_2 output459 (.A(net459),
    .X(soft_irq));
 sky130_fd_sc_hd__buf_2 output460 (.A(net460),
    .X(spim_mosi));
 sky130_fd_sc_hd__buf_2 output461 (.A(net461),
    .X(spis_mosi));
 sky130_fd_sc_hd__buf_2 output462 (.A(net462),
    .X(spis_sck));
 sky130_fd_sc_hd__buf_2 output463 (.A(net463),
    .X(spis_ssn));
 sky130_fd_sc_hd__buf_2 output464 (.A(net464),
    .X(sspim_rst_n));
 sky130_fd_sc_hd__buf_2 output465 (.A(net465),
    .X(strap_sticky[0]));
 sky130_fd_sc_hd__buf_2 output466 (.A(net466),
    .X(strap_sticky[10]));
 sky130_fd_sc_hd__buf_2 output467 (.A(net467),
    .X(strap_sticky[11]));
 sky130_fd_sc_hd__buf_2 output468 (.A(net468),
    .X(strap_sticky[12]));
 sky130_fd_sc_hd__buf_2 output469 (.A(net469),
    .X(strap_sticky[13]));
 sky130_fd_sc_hd__buf_2 output470 (.A(net470),
    .X(strap_sticky[14]));
 sky130_fd_sc_hd__buf_2 output471 (.A(net471),
    .X(strap_sticky[15]));
 sky130_fd_sc_hd__buf_2 output472 (.A(net472),
    .X(strap_sticky[16]));
 sky130_fd_sc_hd__buf_2 output473 (.A(net473),
    .X(strap_sticky[17]));
 sky130_fd_sc_hd__buf_2 output474 (.A(net474),
    .X(strap_sticky[18]));
 sky130_fd_sc_hd__buf_2 output475 (.A(net475),
    .X(strap_sticky[19]));
 sky130_fd_sc_hd__buf_2 output476 (.A(net476),
    .X(strap_sticky[1]));
 sky130_fd_sc_hd__buf_2 output477 (.A(net477),
    .X(strap_sticky[20]));
 sky130_fd_sc_hd__buf_2 output478 (.A(net478),
    .X(strap_sticky[21]));
 sky130_fd_sc_hd__buf_2 output479 (.A(net479),
    .X(strap_sticky[22]));
 sky130_fd_sc_hd__buf_2 output480 (.A(net480),
    .X(strap_sticky[23]));
 sky130_fd_sc_hd__buf_2 output481 (.A(net481),
    .X(strap_sticky[24]));
 sky130_fd_sc_hd__buf_2 output482 (.A(net482),
    .X(strap_sticky[25]));
 sky130_fd_sc_hd__buf_2 output483 (.A(net483),
    .X(strap_sticky[26]));
 sky130_fd_sc_hd__buf_2 output484 (.A(net484),
    .X(strap_sticky[27]));
 sky130_fd_sc_hd__buf_2 output485 (.A(net485),
    .X(strap_sticky[28]));
 sky130_fd_sc_hd__buf_2 output486 (.A(net486),
    .X(strap_sticky[29]));
 sky130_fd_sc_hd__buf_2 output487 (.A(net487),
    .X(strap_sticky[2]));
 sky130_fd_sc_hd__buf_2 output488 (.A(net488),
    .X(strap_sticky[30]));
 sky130_fd_sc_hd__buf_2 output489 (.A(net489),
    .X(strap_sticky[31]));
 sky130_fd_sc_hd__buf_2 output490 (.A(net490),
    .X(strap_sticky[3]));
 sky130_fd_sc_hd__buf_2 output491 (.A(net491),
    .X(strap_sticky[4]));
 sky130_fd_sc_hd__buf_2 output492 (.A(net492),
    .X(strap_sticky[5]));
 sky130_fd_sc_hd__buf_2 output493 (.A(net493),
    .X(strap_sticky[6]));
 sky130_fd_sc_hd__buf_2 output494 (.A(net494),
    .X(strap_sticky[7]));
 sky130_fd_sc_hd__buf_2 output495 (.A(net495),
    .X(strap_sticky[8]));
 sky130_fd_sc_hd__buf_2 output496 (.A(net496),
    .X(strap_sticky[9]));
 sky130_fd_sc_hd__buf_2 output497 (.A(net497),
    .X(strap_uartm[0]));
 sky130_fd_sc_hd__buf_2 output498 (.A(net498),
    .X(strap_uartm[1]));
 sky130_fd_sc_hd__buf_2 output499 (.A(net499),
    .X(uart_rst_n[0]));
 sky130_fd_sc_hd__buf_2 output500 (.A(net500),
    .X(uart_rst_n[1]));
 sky130_fd_sc_hd__buf_2 output501 (.A(net501),
    .X(uart_rxd[0]));
 sky130_fd_sc_hd__buf_2 output502 (.A(net502),
    .X(uart_rxd[1]));
 sky130_fd_sc_hd__buf_2 output503 (.A(net503),
    .X(uartm_rxd));
 sky130_fd_sc_hd__clkbuf_1 output504 (.A(net504),
    .X(usb_clk));
 sky130_fd_sc_hd__buf_2 output505 (.A(net601),
    .X(usb_dn_i));
 sky130_fd_sc_hd__buf_2 output506 (.A(net506),
    .X(usb_dp_i));
 sky130_fd_sc_hd__buf_2 output507 (.A(net507),
    .X(usb_rst_n));
 sky130_fd_sc_hd__buf_2 output508 (.A(net508),
    .X(user_irq[0]));
 sky130_fd_sc_hd__buf_2 output509 (.A(net509),
    .X(user_irq[1]));
 sky130_fd_sc_hd__buf_2 output510 (.A(net510),
    .X(user_irq[2]));
 sky130_fd_sc_hd__buf_2 output511 (.A(net511),
    .X(wbd_clk_pinmux));
 sky130_fd_sc_hd__buf_2 output512 (.A(net512),
    .X(xtal_clk));
 sky130_fd_sc_hd__conb_1 pinmux_top_1657 (.LO(net1657));
 sky130_fd_sc_hd__conb_1 pinmux_top_1658 (.LO(net1658));
 sky130_fd_sc_hd__conb_1 pinmux_top_1659 (.LO(net1659));
 sky130_fd_sc_hd__conb_1 pinmux_top_1660 (.LO(net1660));
 sky130_fd_sc_hd__conb_1 pinmux_top_1661 (.LO(net1661));
 sky130_fd_sc_hd__conb_1 pinmux_top_1662 (.LO(net1662));
 sky130_fd_sc_hd__conb_1 pinmux_top_1663 (.LO(net1663));
 sky130_fd_sc_hd__conb_1 pinmux_top_1664 (.LO(net1664));
 sky130_fd_sc_hd__conb_1 pinmux_top_1665 (.LO(net1665));
 sky130_fd_sc_hd__conb_1 pinmux_top_1666 (.LO(net1666));
 sky130_fd_sc_hd__conb_1 pinmux_top_1667 (.LO(net1667));
 sky130_fd_sc_hd__conb_1 pinmux_top_1668 (.LO(net1668));
 sky130_fd_sc_hd__conb_1 pinmux_top_1669 (.LO(net1669));
 sky130_fd_sc_hd__conb_1 pinmux_top_1670 (.LO(net1670));
 sky130_fd_sc_hd__conb_1 pinmux_top_1671 (.LO(net1671));
 sky130_fd_sc_hd__conb_1 pinmux_top_1672 (.LO(net1672));
 sky130_fd_sc_hd__conb_1 pinmux_top_1673 (.LO(net1673));
 sky130_fd_sc_hd__conb_1 pinmux_top_1674 (.LO(net1674));
 sky130_fd_sc_hd__conb_1 pinmux_top_1675 (.LO(net1675));
 sky130_fd_sc_hd__conb_1 pinmux_top_1676 (.LO(net1676));
 sky130_fd_sc_hd__conb_1 pinmux_top_1677 (.LO(net1677));
 sky130_fd_sc_hd__conb_1 pinmux_top_1678 (.LO(net1678));
 sky130_fd_sc_hd__conb_1 pinmux_top_1679 (.LO(net1679));
 sky130_fd_sc_hd__conb_1 pinmux_top_1680 (.LO(net1680));
 sky130_fd_sc_hd__conb_1 pinmux_top_1681 (.LO(net1681));
 sky130_fd_sc_hd__conb_1 pinmux_top_1682 (.LO(net1682));
 sky130_fd_sc_hd__conb_1 pinmux_top_1683 (.LO(net1683));
 sky130_fd_sc_hd__conb_1 pinmux_top_1684 (.LO(net1684));
 sky130_fd_sc_hd__conb_1 pinmux_top_1685 (.LO(net1685));
 sky130_fd_sc_hd__conb_1 pinmux_top_1686 (.LO(net1686));
 sky130_fd_sc_hd__conb_1 pinmux_top_1687 (.LO(net1687));
 sky130_fd_sc_hd__conb_1 pinmux_top_1688 (.LO(net1688));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer1 (.A(\u_skew_pinmux.clk_d6 ),
    .X(net1700));
 sky130_fd_sc_hd__dlygate4sd1_1 rebuffer2 (.A(\u_skew_pinmux.clk_d7 ),
    .X(net1701));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_cpu0_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[8] ),
    .X(\u_glbl_reg.u_buf_cpu0_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_cpu1_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[9] ),
    .X(\u_glbl_reg.u_buf_cpu1_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_cpu2_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[10] ),
    .X(\u_glbl_reg.u_buf_cpu2_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_cpu3_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[11] ),
    .X(\u_glbl_reg.u_buf_cpu3_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_cpu_intf_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[0] ),
    .X(net252));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_i2cm_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[4] ),
    .X(net331));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_qspim_rst.u_buf  (.A(net1705),
    .X(net367));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_sspim_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[2] ),
    .X(net464));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_uart0_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[3] ),
    .X(\u_glbl_reg.u_buf_uart0_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_uart1_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[6] ),
    .X(\u_glbl_reg.u_buf_uart1_rst.X ));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_buf_usb_rst.u_buf  (.A(\u_glbl_reg.cfg_rst_ctrl[5] ),
    .X(net507));
 sky130_fd_sc_hd__clkbuf_1 \u_glbl_reg.u_clkbuf_dbg.u_buf  (.A(\u_glbl_reg.dbg_clk_div16 ),
    .X(\u_glbl_reg.dbg_clk_mon ));
 sky130_fd_sc_hd__clkbuf_8 \u_glbl_reg.u_clkbuf_dbg_ref.u_buf  (.A(net1693),
    .X(\u_glbl_reg.dbg_clk_ref_buf ));
 sky130_fd_sc_hd__clkbuf_8 \u_glbl_reg.u_clkbuf_rtc.u_buf  (.A(\u_glbl_reg.rtc_clk_int ),
    .X(net454));
 sky130_fd_sc_hd__clkbuf_8 \u_glbl_reg.u_clkbuf_usb.u_buf  (.A(\u_glbl_reg.u_clkbuf_usb.A ),
    .X(net504));
 sky130_fd_sc_hd__mux2_8 \u_glbl_reg.u_rtc_clk_sel.genblk1.u_mux  (.A0(\u_glbl_reg.rtc_ref_clk ),
    .A1(\u_glbl_reg.rtc_clk_div ),
    .S(\u_glbl_reg.cfg_rtc_clk_ctrl[5] ),
    .X(\u_glbl_reg.rtc_clk_int ));
 sky130_fd_sc_hd__clkbuf_8 \u_glbl_reg.u_rtc_ref_clkbuf.u_buf  (.A(\u_glbl_reg.rtc_ref_clk_int ),
    .X(\u_glbl_reg.rtc_ref_clk ));
 sky130_fd_sc_hd__mux2_8 \u_glbl_reg.u_usb_clk_sel.genblk1.u_mux  (.A0(\u_glbl_reg.u_usb_clk_sel.A0 ),
    .A1(\u_glbl_reg.u_usb_clk_sel.A1 ),
    .S(\u_glbl_reg.cfg_usb_clk_ctrl[5] ),
    .X(\u_glbl_reg.u_clkbuf_usb.A ));
 sky130_fd_sc_hd__clkbuf_8 \u_glbl_reg.u_usb_ref_clkbuf.u_buf  (.A(\u_glbl_reg.u_usb_ref_clkbuf.A ),
    .X(\u_glbl_reg.u_usb_clk_sel.A0 ));
 sky130_fd_sc_hd__mux2_1 \u_prst_sync.u_buf.genblk1.u_mux  (.A0(net1843),
    .A1(net48),
    .S(net1655),
    .X(\u_glbl_reg.p_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_prst_sync.u_buf.genblk1.u_mux_1655  (.LO(net1655));
 sky130_fd_sc_hd__mux2_1 \u_rst_sync.u_buf.genblk1.u_mux  (.A0(net1875),
    .A1(net134),
    .S(net1656),
    .X(\u_glbl_reg.s_reset_n ));
 sky130_fd_sc_hd__conb_1 \u_rst_sync.u_buf.genblk1.u_mux_1656  (.LO(net1656));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_1.u_dly0  (.A(\u_skew_pinmux.clk_inbuf ),
    .X(\u_skew_pinmux.clkbuf_1.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_1.u_dly1  (.A(\u_skew_pinmux.clkbuf_1.X1 ),
    .X(\u_skew_pinmux.clkbuf_1.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_1.u_dly2  (.A(\u_skew_pinmux.clkbuf_1.X2 ),
    .X(\u_skew_pinmux.clkbuf_1.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_1.u_dly3  (.A(\u_skew_pinmux.clkbuf_1.X3 ),
    .X(\u_skew_pinmux.clk_d1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_10.u_dly0  (.A(\u_skew_pinmux.clk_d9 ),
    .X(\u_skew_pinmux.clkbuf_10.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_10.u_dly1  (.A(\u_skew_pinmux.clkbuf_10.X1 ),
    .X(\u_skew_pinmux.clkbuf_10.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_10.u_dly2  (.A(\u_skew_pinmux.clkbuf_10.X2 ),
    .X(\u_skew_pinmux.clkbuf_10.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_10.u_dly3  (.A(\u_skew_pinmux.clkbuf_10.X3 ),
    .X(\u_skew_pinmux.clk_d10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_11.u_dly0  (.A(\u_skew_pinmux.clk_d10 ),
    .X(\u_skew_pinmux.clkbuf_11.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_11.u_dly1  (.A(\u_skew_pinmux.clkbuf_11.X1 ),
    .X(\u_skew_pinmux.clkbuf_11.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_11.u_dly2  (.A(\u_skew_pinmux.clkbuf_11.X2 ),
    .X(\u_skew_pinmux.clkbuf_11.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_11.u_dly3  (.A(\u_skew_pinmux.clkbuf_11.X3 ),
    .X(\u_skew_pinmux.clk_d11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_12.u_dly0  (.A(\u_skew_pinmux.clk_d11 ),
    .X(\u_skew_pinmux.clkbuf_12.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_12.u_dly1  (.A(\u_skew_pinmux.clkbuf_12.X1 ),
    .X(\u_skew_pinmux.clkbuf_12.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_12.u_dly2  (.A(\u_skew_pinmux.clkbuf_12.X2 ),
    .X(\u_skew_pinmux.clkbuf_12.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_12.u_dly3  (.A(\u_skew_pinmux.clkbuf_12.X3 ),
    .X(\u_skew_pinmux.clk_d12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_13.u_dly0  (.A(\u_skew_pinmux.clk_d12 ),
    .X(\u_skew_pinmux.clkbuf_13.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_13.u_dly1  (.A(\u_skew_pinmux.clkbuf_13.X1 ),
    .X(\u_skew_pinmux.clkbuf_13.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_13.u_dly2  (.A(\u_skew_pinmux.clkbuf_13.X2 ),
    .X(\u_skew_pinmux.clkbuf_13.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_13.u_dly3  (.A(\u_skew_pinmux.clkbuf_13.X3 ),
    .X(\u_skew_pinmux.clk_d13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_14.u_dly0  (.A(\u_skew_pinmux.clk_d13 ),
    .X(\u_skew_pinmux.clkbuf_14.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_14.u_dly1  (.A(\u_skew_pinmux.clkbuf_14.X1 ),
    .X(\u_skew_pinmux.clkbuf_14.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_14.u_dly2  (.A(\u_skew_pinmux.clkbuf_14.X2 ),
    .X(\u_skew_pinmux.clkbuf_14.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_14.u_dly3  (.A(\u_skew_pinmux.clkbuf_14.X3 ),
    .X(\u_skew_pinmux.clk_d14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_15.u_dly0  (.A(\u_skew_pinmux.clk_d14 ),
    .X(\u_skew_pinmux.clkbuf_15.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_15.u_dly1  (.A(\u_skew_pinmux.clkbuf_15.X1 ),
    .X(\u_skew_pinmux.clkbuf_15.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_15.u_dly2  (.A(\u_skew_pinmux.clkbuf_15.X2 ),
    .X(\u_skew_pinmux.clkbuf_15.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_15.u_dly3  (.A(\u_skew_pinmux.clkbuf_15.X3 ),
    .X(\u_skew_pinmux.clk_d15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_2.u_dly0  (.A(\u_skew_pinmux.clk_d1 ),
    .X(\u_skew_pinmux.clkbuf_2.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_2.u_dly1  (.A(\u_skew_pinmux.clkbuf_2.X1 ),
    .X(\u_skew_pinmux.clkbuf_2.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_2.u_dly2  (.A(\u_skew_pinmux.clkbuf_2.X2 ),
    .X(\u_skew_pinmux.clkbuf_2.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_2.u_dly3  (.A(\u_skew_pinmux.clkbuf_2.X3 ),
    .X(\u_skew_pinmux.clk_d2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_3.u_dly0  (.A(\u_skew_pinmux.clk_d2 ),
    .X(\u_skew_pinmux.clkbuf_3.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_3.u_dly1  (.A(\u_skew_pinmux.clkbuf_3.X1 ),
    .X(\u_skew_pinmux.clkbuf_3.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_3.u_dly2  (.A(\u_skew_pinmux.clkbuf_3.X2 ),
    .X(\u_skew_pinmux.clkbuf_3.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_3.u_dly3  (.A(\u_skew_pinmux.clkbuf_3.X3 ),
    .X(\u_skew_pinmux.clk_d3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_4.u_dly0  (.A(\u_skew_pinmux.clk_d3 ),
    .X(\u_skew_pinmux.clkbuf_4.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_4.u_dly1  (.A(\u_skew_pinmux.clkbuf_4.X1 ),
    .X(\u_skew_pinmux.clkbuf_4.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_4.u_dly2  (.A(\u_skew_pinmux.clkbuf_4.X2 ),
    .X(\u_skew_pinmux.clkbuf_4.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_4.u_dly3  (.A(\u_skew_pinmux.clkbuf_4.X3 ),
    .X(\u_skew_pinmux.clk_d4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_5.u_dly0  (.A(\u_skew_pinmux.clk_d4 ),
    .X(\u_skew_pinmux.clkbuf_5.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_5.u_dly1  (.A(\u_skew_pinmux.clkbuf_5.X1 ),
    .X(\u_skew_pinmux.clkbuf_5.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_5.u_dly2  (.A(\u_skew_pinmux.clkbuf_5.X2 ),
    .X(\u_skew_pinmux.clkbuf_5.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_5.u_dly3  (.A(\u_skew_pinmux.clkbuf_5.X3 ),
    .X(\u_skew_pinmux.clk_d5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_6.u_dly0  (.A(\u_skew_pinmux.clk_d5 ),
    .X(\u_skew_pinmux.clkbuf_6.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_6.u_dly1  (.A(\u_skew_pinmux.clkbuf_6.X1 ),
    .X(\u_skew_pinmux.clkbuf_6.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_6.u_dly2  (.A(\u_skew_pinmux.clkbuf_6.X2 ),
    .X(\u_skew_pinmux.clkbuf_6.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_6.u_dly3  (.A(\u_skew_pinmux.clkbuf_6.X3 ),
    .X(\u_skew_pinmux.clk_d6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_7.u_dly0  (.A(\u_skew_pinmux.clk_d6 ),
    .X(\u_skew_pinmux.clkbuf_7.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_7.u_dly1  (.A(\u_skew_pinmux.clkbuf_7.X1 ),
    .X(\u_skew_pinmux.clkbuf_7.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_7.u_dly2  (.A(\u_skew_pinmux.clkbuf_7.X2 ),
    .X(\u_skew_pinmux.clkbuf_7.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_7.u_dly3  (.A(\u_skew_pinmux.clkbuf_7.X3 ),
    .X(\u_skew_pinmux.clk_d7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_8.u_dly0  (.A(\u_skew_pinmux.clk_d7 ),
    .X(\u_skew_pinmux.clkbuf_8.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_8.u_dly1  (.A(\u_skew_pinmux.clkbuf_8.X1 ),
    .X(\u_skew_pinmux.clkbuf_8.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_8.u_dly2  (.A(\u_skew_pinmux.clkbuf_8.X2 ),
    .X(\u_skew_pinmux.clkbuf_8.X3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_8.u_dly3  (.A(\u_skew_pinmux.clkbuf_8.X3 ),
    .X(\u_skew_pinmux.clk_d8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_9.u_dly0  (.A(\u_skew_pinmux.clk_d8 ),
    .X(\u_skew_pinmux.clkbuf_9.X1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_9.u_dly1  (.A(\u_skew_pinmux.clkbuf_9.X1 ),
    .X(\u_skew_pinmux.clkbuf_9.X2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.clkbuf_9.u_dly2  (.A(\u_skew_pinmux.clkbuf_9.X2 ),
    .X(\u_skew_pinmux.clkbuf_9.X3 ));
 sky130_fd_sc_hd__buf_2 \u_skew_pinmux.clkbuf_9.u_dly3  (.A(\u_skew_pinmux.clkbuf_9.X3 ),
    .X(\u_skew_pinmux.clk_d9 ));
 sky130_fd_sc_hd__buf_6 \u_skew_pinmux.u_clkbuf_in.u_buf  (.A(net198),
    .X(\u_skew_pinmux.clk_inbuf ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_clkbuf_out.u_buf  (.A(\u_skew_pinmux.d30 ),
    .X(net511));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_00.genblk1.u_mux  (.A0(\u_skew_pinmux.in0 ),
    .A1(\u_skew_pinmux.in1 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d00 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_01.genblk1.u_mux  (.A0(\u_skew_pinmux.in2 ),
    .A1(\u_skew_pinmux.in3 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d01 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_02.genblk1.u_mux  (.A0(\u_skew_pinmux.in4 ),
    .A1(\u_skew_pinmux.in5 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d02 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_03.genblk1.u_mux  (.A0(\u_skew_pinmux.in6 ),
    .A1(\u_skew_pinmux.in7 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d03 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_04.genblk1.u_mux  (.A0(\u_skew_pinmux.in8 ),
    .A1(\u_skew_pinmux.in9 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d04 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_05.genblk1.u_mux  (.A0(\u_skew_pinmux.in10 ),
    .A1(\u_skew_pinmux.in11 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d05 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_06.genblk1.u_mux  (.A0(\u_skew_pinmux.in12 ),
    .A1(\u_skew_pinmux.in13 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d06 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_07.genblk1.u_mux  (.A0(\u_skew_pinmux.in14 ),
    .A1(\u_skew_pinmux.in15 ),
    .S(cfg_cska_pinmux[0]),
    .X(\u_skew_pinmux.d07 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_10.genblk1.u_mux  (.A0(\u_skew_pinmux.d00 ),
    .A1(\u_skew_pinmux.d01 ),
    .S(cfg_cska_pinmux[1]),
    .X(\u_skew_pinmux.d10 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_11.genblk1.u_mux  (.A0(\u_skew_pinmux.d02 ),
    .A1(\u_skew_pinmux.d03 ),
    .S(cfg_cska_pinmux[1]),
    .X(\u_skew_pinmux.d11 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_12.genblk1.u_mux  (.A0(\u_skew_pinmux.d04 ),
    .A1(\u_skew_pinmux.d05 ),
    .S(cfg_cska_pinmux[1]),
    .X(\u_skew_pinmux.d12 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_13.genblk1.u_mux  (.A0(\u_skew_pinmux.d06 ),
    .A1(\u_skew_pinmux.d07 ),
    .S(cfg_cska_pinmux[1]),
    .X(\u_skew_pinmux.d13 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_20.genblk1.u_mux  (.A0(\u_skew_pinmux.d10 ),
    .A1(\u_skew_pinmux.d11 ),
    .S(cfg_cska_pinmux[2]),
    .X(\u_skew_pinmux.d20 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_21.genblk1.u_mux  (.A0(\u_skew_pinmux.d12 ),
    .A1(\u_skew_pinmux.d13 ),
    .S(cfg_cska_pinmux[2]),
    .X(\u_skew_pinmux.d21 ));
 sky130_fd_sc_hd__mux2_1 \u_skew_pinmux.u_mux_level_30.genblk1.u_mux  (.A0(\u_skew_pinmux.d20 ),
    .A1(\u_skew_pinmux.d21 ),
    .S(cfg_cska_pinmux[3]),
    .X(\u_skew_pinmux.d30 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_0.u_buf  (.A(\u_skew_pinmux.clk_inbuf ),
    .X(\u_skew_pinmux.in0 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_1.u_buf  (.A(\u_skew_pinmux.clk_d1 ),
    .X(\u_skew_pinmux.in1 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_10.u_buf  (.A(\u_skew_pinmux.clk_d10 ),
    .X(\u_skew_pinmux.in10 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_11.u_buf  (.A(\u_skew_pinmux.clk_d11 ),
    .X(\u_skew_pinmux.in11 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_12.u_buf  (.A(\u_skew_pinmux.clk_d12 ),
    .X(\u_skew_pinmux.in12 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_13.u_buf  (.A(\u_skew_pinmux.clk_d13 ),
    .X(\u_skew_pinmux.in13 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_14.u_buf  (.A(\u_skew_pinmux.clk_d14 ),
    .X(\u_skew_pinmux.in14 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_15.u_buf  (.A(\u_skew_pinmux.clk_d15 ),
    .X(\u_skew_pinmux.in15 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_2.u_buf  (.A(\u_skew_pinmux.clk_d2 ),
    .X(\u_skew_pinmux.in2 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_3.u_buf  (.A(\u_skew_pinmux.clk_d3 ),
    .X(\u_skew_pinmux.in3 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_4.u_buf  (.A(\u_skew_pinmux.clk_d4 ),
    .X(\u_skew_pinmux.in4 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_5.u_buf  (.A(\u_skew_pinmux.clk_d5 ),
    .X(\u_skew_pinmux.in5 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_6.u_buf  (.A(net1700),
    .X(\u_skew_pinmux.in6 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_7.u_buf  (.A(net1701),
    .X(\u_skew_pinmux.in7 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_8.u_buf  (.A(\u_skew_pinmux.clk_d8 ),
    .X(\u_skew_pinmux.in8 ));
 sky130_fd_sc_hd__clkbuf_1 \u_skew_pinmux.u_tap_9.u_buf  (.A(\u_skew_pinmux.clk_d9 ),
    .X(\u_skew_pinmux.in9 ));
 sky130_fd_sc_hd__buf_4 wire1043 (.A(net1042),
    .X(net1043));
 sky130_fd_sc_hd__buf_6 wire1069 (.A(net1068),
    .X(net1069));
 sky130_fd_sc_hd__buf_6 wire1078 (.A(\u_ws281x.u_txd_1.txd ),
    .X(net1078));
 sky130_fd_sc_hd__buf_6 wire1079 (.A(\u_ws281x.u_txd_0.txd ),
    .X(net1079));
 sky130_fd_sc_hd__buf_4 wire1093 (.A(net222),
    .X(net1093));
 sky130_fd_sc_hd__buf_4 wire1094 (.A(net221),
    .X(net1094));
 sky130_fd_sc_hd__buf_4 wire1095 (.A(net220),
    .X(net1095));
 sky130_fd_sc_hd__buf_4 wire1096 (.A(net219),
    .X(net1096));
 sky130_fd_sc_hd__buf_4 wire1097 (.A(net218),
    .X(net1097));
 sky130_fd_sc_hd__clkbuf_4 wire1098 (.A(net217),
    .X(net1098));
 sky130_fd_sc_hd__buf_4 wire1099 (.A(net210),
    .X(net1099));
 sky130_fd_sc_hd__buf_4 wire1100 (.A(net225),
    .X(net1100));
 sky130_fd_sc_hd__buf_4 wire1101 (.A(net231),
    .X(net1101));
 sky130_fd_sc_hd__buf_4 wire1102 (.A(net230),
    .X(net1102));
 sky130_fd_sc_hd__buf_4 wire1103 (.A(net229),
    .X(net1103));
 sky130_fd_sc_hd__buf_4 wire1104 (.A(net228),
    .X(net1104));
 sky130_fd_sc_hd__buf_4 wire1105 (.A(net227),
    .X(net1105));
 sky130_fd_sc_hd__buf_4 wire1106 (.A(net216),
    .X(net1106));
 sky130_fd_sc_hd__buf_4 wire1107 (.A(net215),
    .X(net1107));
 sky130_fd_sc_hd__buf_4 wire1108 (.A(net226),
    .X(net1108));
 sky130_fd_sc_hd__buf_6 wire1183 (.A(net1184),
    .X(net1183));
 sky130_fd_sc_hd__buf_6 wire1184 (.A(net320),
    .X(net1184));
 sky130_fd_sc_hd__buf_6 wire1185 (.A(net1186),
    .X(net1185));
 sky130_fd_sc_hd__buf_6 wire1186 (.A(net319),
    .X(net1186));
 sky130_fd_sc_hd__buf_6 wire1187 (.A(net1188),
    .X(net1187));
 sky130_fd_sc_hd__buf_6 wire1188 (.A(net318),
    .X(net1188));
 sky130_fd_sc_hd__buf_6 wire1189 (.A(net1190),
    .X(net1189));
 sky130_fd_sc_hd__buf_6 wire1190 (.A(net317),
    .X(net1190));
 sky130_fd_sc_hd__buf_6 wire1191 (.A(net1192),
    .X(net1191));
 sky130_fd_sc_hd__buf_6 wire1192 (.A(net316),
    .X(net1192));
 sky130_fd_sc_hd__buf_6 wire1193 (.A(net1194),
    .X(net1193));
 sky130_fd_sc_hd__buf_6 wire1194 (.A(net315),
    .X(net1194));
 sky130_fd_sc_hd__buf_6 wire1195 (.A(net1196),
    .X(net1195));
 sky130_fd_sc_hd__buf_6 wire1196 (.A(net314),
    .X(net1196));
 sky130_fd_sc_hd__buf_6 wire1197 (.A(net1198),
    .X(net1197));
 sky130_fd_sc_hd__buf_6 wire1198 (.A(net312),
    .X(net1198));
 sky130_fd_sc_hd__buf_6 wire1199 (.A(net1200),
    .X(net1199));
 sky130_fd_sc_hd__buf_6 wire1200 (.A(net311),
    .X(net1200));
 sky130_fd_sc_hd__buf_6 wire1206 (.A(net365),
    .X(net1206));
 sky130_fd_sc_hd__buf_4 wire1285 (.A(net1284),
    .X(net1285));
 sky130_fd_sc_hd__buf_4 wire1292 (.A(net99),
    .X(net1292));
 sky130_fd_sc_hd__buf_6 wire1304 (.A(net9),
    .X(net1304));
 sky130_fd_sc_hd__buf_4 wire1305 (.A(net8),
    .X(net1305));
 sky130_fd_sc_hd__buf_4 wire1306 (.A(net7),
    .X(net1306));
 sky130_fd_sc_hd__buf_6 wire1307 (.A(net64),
    .X(net1307));
 sky130_fd_sc_hd__buf_4 wire1314 (.A(net1312),
    .X(net1314));
 sky130_fd_sc_hd__buf_4 wire1315 (.A(net63),
    .X(net1315));
 sky130_fd_sc_hd__buf_6 wire1318 (.A(net1317),
    .X(net1318));
 sky130_fd_sc_hd__buf_4 wire1327 (.A(net1326),
    .X(net1327));
 sky130_fd_sc_hd__clkbuf_8 wire1330 (.A(net61),
    .X(net1330));
 sky130_fd_sc_hd__buf_4 wire1338 (.A(net60),
    .X(net1338));
 sky130_fd_sc_hd__buf_6 wire1339 (.A(net6),
    .X(net1339));
 sky130_fd_sc_hd__buf_6 wire1340 (.A(net59),
    .X(net1340));
 sky130_fd_sc_hd__buf_6 wire1341 (.A(net58),
    .X(net1341));
 sky130_fd_sc_hd__buf_8 wire1342 (.A(net57),
    .X(net1342));
 sky130_fd_sc_hd__buf_6 wire1345 (.A(net55),
    .X(net1345));
 sky130_fd_sc_hd__buf_4 wire1347 (.A(net54),
    .X(net1347));
 sky130_fd_sc_hd__clkbuf_4 wire1373 (.A(net51),
    .X(net1373));
 sky130_fd_sc_hd__buf_6 wire1374 (.A(net50),
    .X(net1374));
 sky130_fd_sc_hd__buf_6 wire1375 (.A(net5),
    .X(net1375));
 sky130_fd_sc_hd__clkbuf_4 wire1376 (.A(net49),
    .X(net1376));
 sky130_fd_sc_hd__clkbuf_4 wire1377 (.A(net40),
    .X(net1377));
 sky130_fd_sc_hd__buf_8 wire1386 (.A(net1385),
    .X(net1386));
 sky130_fd_sc_hd__buf_4 wire1387 (.A(net37),
    .X(net1387));
 sky130_fd_sc_hd__buf_6 wire1388 (.A(net35),
    .X(net1388));
 sky130_fd_sc_hd__buf_4 wire1389 (.A(net1390),
    .X(net1389));
 sky130_fd_sc_hd__buf_6 wire1390 (.A(net31),
    .X(net1390));
 sky130_fd_sc_hd__buf_6 wire1391 (.A(net30),
    .X(net1391));
 sky130_fd_sc_hd__buf_4 wire1392 (.A(net3),
    .X(net1392));
 sky130_fd_sc_hd__buf_4 wire1393 (.A(net1394),
    .X(net1393));
 sky130_fd_sc_hd__buf_6 wire1394 (.A(net29),
    .X(net1394));
 sky130_fd_sc_hd__buf_4 wire1395 (.A(net1396),
    .X(net1395));
 sky130_fd_sc_hd__buf_6 wire1396 (.A(net28),
    .X(net1396));
 sky130_fd_sc_hd__clkbuf_4 wire1397 (.A(net23),
    .X(net1397));
 sky130_fd_sc_hd__clkbuf_4 wire1398 (.A(net197),
    .X(net1398));
 sky130_fd_sc_hd__clkbuf_4 wire1399 (.A(net194),
    .X(net1399));
 sky130_fd_sc_hd__buf_8 wire1400 (.A(net16),
    .X(net1400));
 sky130_fd_sc_hd__buf_4 wire1401 (.A(net151),
    .X(net1401));
 sky130_fd_sc_hd__buf_4 wire1402 (.A(net150),
    .X(net1402));
 sky130_fd_sc_hd__buf_8 wire1403 (.A(net15),
    .X(net1403));
 sky130_fd_sc_hd__buf_4 wire1404 (.A(net149),
    .X(net1404));
 sky130_fd_sc_hd__buf_4 wire1405 (.A(net148),
    .X(net1405));
 sky130_fd_sc_hd__buf_6 wire1406 (.A(net1407),
    .X(net1406));
 sky130_fd_sc_hd__buf_6 wire1407 (.A(net142),
    .X(net1407));
 sky130_fd_sc_hd__buf_6 wire1408 (.A(net1409),
    .X(net1408));
 sky130_fd_sc_hd__buf_6 wire1409 (.A(net141),
    .X(net1409));
 sky130_fd_sc_hd__buf_6 wire1410 (.A(net1411),
    .X(net1410));
 sky130_fd_sc_hd__buf_6 wire1411 (.A(net140),
    .X(net1411));
 sky130_fd_sc_hd__buf_6 wire1412 (.A(net1413),
    .X(net1412));
 sky130_fd_sc_hd__buf_6 wire1413 (.A(net139),
    .X(net1413));
 sky130_fd_sc_hd__buf_4 wire1414 (.A(net132),
    .X(net1414));
 sky130_fd_sc_hd__buf_4 wire1415 (.A(net131),
    .X(net1415));
 sky130_fd_sc_hd__buf_4 wire1416 (.A(net130),
    .X(net1416));
 sky130_fd_sc_hd__buf_6 wire1417 (.A(net13),
    .X(net1417));
 sky130_fd_sc_hd__buf_4 wire1424 (.A(net129),
    .X(net1424));
 sky130_fd_sc_hd__buf_4 wire1432 (.A(net1430),
    .X(net1432));
 sky130_fd_sc_hd__buf_4 wire1439 (.A(net1438),
    .X(net1439));
 sky130_fd_sc_hd__buf_4 wire1455 (.A(net1454),
    .X(net1455));
 sky130_fd_sc_hd__buf_4 wire1456 (.A(net125),
    .X(net1456));
 sky130_fd_sc_hd__buf_4 wire1464 (.A(net1463),
    .X(net1464));
 sky130_fd_sc_hd__buf_4 wire1465 (.A(net124),
    .X(net1465));
 sky130_fd_sc_hd__buf_6 wire1472 (.A(net1471),
    .X(net1472));
 sky130_fd_sc_hd__buf_4 wire1473 (.A(net123),
    .X(net1473));
 sky130_fd_sc_hd__buf_6 wire1480 (.A(net1479),
    .X(net1480));
 sky130_fd_sc_hd__buf_8 wire1487 (.A(net1486),
    .X(net1487));
 sky130_fd_sc_hd__buf_4 wire1495 (.A(net1494),
    .X(net1495));
 sky130_fd_sc_hd__buf_6 wire1497 (.A(net12),
    .X(net1497));
 sky130_fd_sc_hd__buf_8 wire1504 (.A(net1503),
    .X(net1504));
 sky130_fd_sc_hd__buf_8 wire1511 (.A(net1510),
    .X(net1511));
 sky130_fd_sc_hd__buf_6 wire1518 (.A(net1517),
    .X(net1518));
 sky130_fd_sc_hd__buf_6 wire1525 (.A(net1524),
    .X(net1525));
 sky130_fd_sc_hd__buf_4 wire1532 (.A(net1533),
    .X(net1532));
 sky130_fd_sc_hd__buf_4 wire1533 (.A(net1531),
    .X(net1533));
 sky130_fd_sc_hd__buf_8 wire1540 (.A(net1539),
    .X(net1540));
 sky130_fd_sc_hd__buf_4 wire1544 (.A(net1543),
    .X(net1544));
 sky130_fd_sc_hd__buf_4 wire1563 (.A(net1562),
    .X(net1563));
 sky130_fd_sc_hd__buf_6 wire1571 (.A(net11),
    .X(net1571));
 sky130_fd_sc_hd__buf_4 wire1578 (.A(net1577),
    .X(net1578));
 sky130_fd_sc_hd__clkbuf_8 wire1585 (.A(net1584),
    .X(net1585));
 sky130_fd_sc_hd__buf_4 wire1588 (.A(net1587),
    .X(net1588));
 sky130_fd_sc_hd__buf_4 wire1593 (.A(net1592),
    .X(net1593));
 sky130_fd_sc_hd__buf_4 wire1594 (.A(net107),
    .X(net1594));
 sky130_fd_sc_hd__buf_4 wire1596 (.A(net1595),
    .X(net1596));
 sky130_fd_sc_hd__buf_6 wire1605 (.A(net1604),
    .X(net1605));
 sky130_fd_sc_hd__buf_4 wire1609 (.A(net1608),
    .X(net1609));
 sky130_fd_sc_hd__buf_4 wire1611 (.A(net1610),
    .X(net1611));
 sky130_fd_sc_hd__clkbuf_4 wire1612 (.A(net1610),
    .X(net1612));
 sky130_fd_sc_hd__buf_6 wire1620 (.A(net1619),
    .X(net1620));
 sky130_fd_sc_hd__buf_4 wire1627 (.A(net1626),
    .X(net1627));
 sky130_fd_sc_hd__buf_4 wire1634 (.A(net1635),
    .X(net1634));
 sky130_fd_sc_hd__buf_4 wire1635 (.A(net1633),
    .X(net1635));
 sky130_fd_sc_hd__buf_4 wire1642 (.A(net1641),
    .X(net1642));
 sky130_fd_sc_hd__buf_4 wire1649 (.A(net1648),
    .X(net1649));
 sky130_fd_sc_hd__buf_6 wire1650 (.A(net10),
    .X(net1650));
 sky130_fd_sc_hd__buf_4 wire1652 (.A(net1651),
    .X(net1652));
 sky130_fd_sc_hd__buf_4 wire1653 (.A(net1),
    .X(net1653));
 sky130_fd_sc_hd__buf_2 wire2 (.A(mclk),
    .X(net1692));
 sky130_fd_sc_hd__buf_4 wire3 (.A(net1694),
    .X(net1693));
 sky130_fd_sc_hd__clkbuf_2 wire4 (.A(\u_glbl_reg.dbg_clk_ref ),
    .X(net1694));
 sky130_fd_sc_hd__buf_4 wire527 (.A(net301),
    .X(net527));
 sky130_fd_sc_hd__buf_4 wire528 (.A(net326),
    .X(net528));
 sky130_fd_sc_hd__clkbuf_4 wire529 (.A(net296),
    .X(net529));
 sky130_fd_sc_hd__buf_4 wire530 (.A(net299),
    .X(net530));
 sky130_fd_sc_hd__buf_4 wire531 (.A(net300),
    .X(net531));
 sky130_fd_sc_hd__buf_4 wire532 (.A(net303),
    .X(net532));
 sky130_fd_sc_hd__buf_4 wire533 (.A(net366),
    .X(net533));
 sky130_fd_sc_hd__buf_4 wire536 (.A(net261),
    .X(net536));
 sky130_fd_sc_hd__buf_4 wire537 (.A(net262),
    .X(net537));
 sky130_fd_sc_hd__buf_4 wire538 (.A(net263),
    .X(net538));
 sky130_fd_sc_hd__clkbuf_4 wire564 (.A(_01594_),
    .X(net564));
 sky130_fd_sc_hd__buf_4 wire565 (.A(net298),
    .X(net565));
 sky130_fd_sc_hd__buf_4 wire566 (.A(net304),
    .X(net566));
 sky130_fd_sc_hd__buf_4 wire567 (.A(_01340_),
    .X(net567));
 sky130_fd_sc_hd__buf_4 wire581 (.A(net259),
    .X(net581));
 sky130_fd_sc_hd__buf_4 wire582 (.A(net260),
    .X(net582));
 sky130_fd_sc_hd__buf_4 wire583 (.A(net265),
    .X(net583));
 sky130_fd_sc_hd__clkbuf_4 wire6 (.A(clknet_0_mclk),
    .X(net1696));
 sky130_fd_sc_hd__clkbuf_4 wire601 (.A(net505),
    .X(net601));
 sky130_fd_sc_hd__buf_4 wire602 (.A(net266),
    .X(net602));
 sky130_fd_sc_hd__buf_4 wire7 (.A(net1698),
    .X(net1697));
 sky130_fd_sc_hd__clkbuf_2 wire8 (.A(net1699),
    .X(net1698));
 sky130_fd_sc_hd__clkbuf_2 wire9 (.A(net454),
    .X(net1699));
 assign pinmux_debug[0] = net1657;
 assign pinmux_debug[10] = net1667;
 assign pinmux_debug[11] = net1668;
 assign pinmux_debug[12] = net1669;
 assign pinmux_debug[13] = net1670;
 assign pinmux_debug[14] = net1671;
 assign pinmux_debug[15] = net1672;
 assign pinmux_debug[16] = net1673;
 assign pinmux_debug[17] = net1674;
 assign pinmux_debug[18] = net1675;
 assign pinmux_debug[19] = net1676;
 assign pinmux_debug[1] = net1658;
 assign pinmux_debug[20] = net1677;
 assign pinmux_debug[21] = net1678;
 assign pinmux_debug[22] = net1679;
 assign pinmux_debug[23] = net1680;
 assign pinmux_debug[24] = net1681;
 assign pinmux_debug[25] = net1682;
 assign pinmux_debug[26] = net1683;
 assign pinmux_debug[27] = net1684;
 assign pinmux_debug[28] = net1685;
 assign pinmux_debug[29] = net1686;
 assign pinmux_debug[2] = net1659;
 assign pinmux_debug[30] = net1687;
 assign pinmux_debug[31] = net1688;
 assign pinmux_debug[3] = net1660;
 assign pinmux_debug[4] = net1661;
 assign pinmux_debug[5] = net1662;
 assign pinmux_debug[6] = net1663;
 assign pinmux_debug[7] = net1664;
 assign pinmux_debug[8] = net1665;
 assign pinmux_debug[9] = net1666;
endmodule

