magic
tech sky130A
magscale 1 2
timestamp 1698759052
<< obsli1 >>
rect 1104 2159 102856 157777
<< obsm1 >>
rect 14 8 103118 159588
<< metal2 >>
rect 110 159200 166 160800
rect 294 159200 350 160800
rect 478 159200 534 160800
rect 662 159200 718 160800
rect 846 159200 902 160800
rect 1030 159200 1086 160800
rect 1214 159200 1270 160800
rect 1398 159200 1454 160800
rect 1582 159200 1638 160800
rect 1766 159200 1822 160800
rect 1950 159200 2006 160800
rect 2134 159200 2190 160800
rect 2318 159200 2374 160800
rect 2502 159200 2558 160800
rect 2686 159200 2742 160800
rect 2870 159200 2926 160800
rect 3054 159200 3110 160800
rect 3238 159200 3294 160800
rect 3422 159200 3478 160800
rect 3606 159200 3662 160800
rect 3790 159200 3846 160800
rect 3974 159200 4030 160800
rect 4158 159200 4214 160800
rect 4342 159200 4398 160800
rect 4526 159200 4582 160800
rect 4710 159200 4766 160800
rect 4894 159200 4950 160800
rect 5078 159200 5134 160800
rect 5262 159200 5318 160800
rect 5446 159200 5502 160800
rect 5630 159200 5686 160800
rect 5814 159200 5870 160800
rect 5998 159200 6054 160800
rect 6182 159200 6238 160800
rect 6366 159200 6422 160800
rect 6550 159200 6606 160800
rect 6734 159200 6790 160800
rect 6918 159200 6974 160800
rect 7102 159200 7158 160800
rect 7286 159200 7342 160800
rect 7470 159200 7526 160800
rect 7654 159200 7710 160800
rect 30102 159200 30158 160800
rect 30286 159200 30342 160800
rect 30470 159200 30526 160800
rect 30654 159200 30710 160800
rect 30838 159200 30894 160800
rect 31022 159200 31078 160800
rect 31206 159200 31262 160800
rect 31390 159200 31446 160800
rect 31574 159200 31630 160800
rect 40038 159200 40094 160800
rect 40222 159200 40278 160800
rect 40406 159200 40462 160800
rect 40590 159200 40646 160800
rect 40774 159200 40830 160800
rect 40958 159200 41014 160800
rect 41142 159200 41198 160800
rect 41326 159200 41382 160800
rect 41510 159200 41566 160800
rect 41694 159200 41750 160800
rect 41878 159200 41934 160800
rect 42062 159200 42118 160800
rect 42246 159200 42302 160800
rect 42430 159200 42486 160800
rect 42614 159200 42670 160800
rect 42798 159200 42854 160800
rect 42982 159200 43038 160800
rect 43166 159200 43222 160800
rect 43350 159200 43406 160800
rect 43534 159200 43590 160800
rect 43718 159200 43774 160800
rect 43902 159200 43958 160800
rect 44086 159200 44142 160800
rect 44270 159200 44326 160800
rect 44454 159200 44510 160800
rect 44638 159200 44694 160800
rect 44822 159200 44878 160800
rect 45006 159200 45062 160800
rect 45190 159200 45246 160800
rect 45374 159200 45430 160800
rect 45558 159200 45614 160800
rect 45742 159200 45798 160800
rect 45926 159200 45982 160800
rect 46110 159200 46166 160800
rect 46294 159200 46350 160800
rect 46478 159200 46534 160800
rect 46662 159200 46718 160800
rect 46846 159200 46902 160800
rect 47030 159200 47086 160800
rect 47214 159200 47270 160800
rect 47398 159200 47454 160800
rect 47582 159200 47638 160800
rect 47766 159200 47822 160800
rect 47950 159200 48006 160800
rect 48134 159200 48190 160800
rect 48318 159200 48374 160800
rect 48502 159200 48558 160800
rect 48686 159200 48742 160800
rect 48870 159200 48926 160800
rect 49054 159200 49110 160800
rect 49238 159200 49294 160800
rect 49422 159200 49478 160800
rect 49606 159200 49662 160800
rect 49790 159200 49846 160800
rect 49974 159200 50030 160800
rect 50158 159200 50214 160800
rect 50342 159200 50398 160800
rect 50526 159200 50582 160800
rect 50710 159200 50766 160800
rect 50894 159200 50950 160800
rect 51078 159200 51134 160800
rect 51262 159200 51318 160800
rect 51446 159200 51502 160800
rect 51630 159200 51686 160800
rect 51814 159200 51870 160800
rect 51998 159200 52054 160800
rect 52182 159200 52238 160800
rect 52366 159200 52422 160800
rect 52550 159200 52606 160800
rect 52734 159200 52790 160800
rect 52918 159200 52974 160800
rect 53102 159200 53158 160800
rect 53286 159200 53342 160800
rect 53470 159200 53526 160800
rect 53654 159200 53710 160800
rect 53838 159200 53894 160800
rect 54022 159200 54078 160800
rect 54206 159200 54262 160800
rect 54390 159200 54446 160800
rect 54574 159200 54630 160800
rect 54758 159200 54814 160800
rect 54942 159200 54998 160800
rect 60094 159200 60150 160800
rect 60278 159200 60334 160800
rect 60462 159200 60518 160800
rect 60646 159200 60702 160800
rect 60830 159200 60886 160800
rect 61014 159200 61070 160800
rect 61198 159200 61254 160800
rect 61382 159200 61438 160800
rect 61566 159200 61622 160800
rect 61750 159200 61806 160800
rect 61934 159200 61990 160800
rect 62118 159200 62174 160800
rect 62302 159200 62358 160800
rect 62486 159200 62542 160800
rect 62670 159200 62726 160800
rect 62854 159200 62910 160800
rect 63038 159200 63094 160800
rect 63222 159200 63278 160800
rect 63406 159200 63462 160800
rect 63590 159200 63646 160800
rect 63774 159200 63830 160800
rect 63958 159200 64014 160800
rect 64142 159200 64198 160800
rect 64326 159200 64382 160800
rect 64510 159200 64566 160800
rect 64694 159200 64750 160800
rect 64878 159200 64934 160800
rect 65062 159200 65118 160800
rect 65246 159200 65302 160800
rect 65430 159200 65486 160800
rect 65614 159200 65670 160800
rect 65798 159200 65854 160800
rect 65982 159200 66038 160800
rect 66166 159200 66222 160800
rect 80058 159200 80114 160800
rect 80242 159200 80298 160800
rect 80426 159200 80482 160800
rect 80610 159200 80666 160800
rect 80794 159200 80850 160800
rect 80978 159200 81034 160800
rect 81162 159200 81218 160800
rect 81346 159200 81402 160800
rect 81530 159200 81586 160800
rect 81714 159200 81770 160800
rect 81898 159200 81954 160800
rect 82082 159200 82138 160800
rect 82266 159200 82322 160800
rect 82450 159200 82506 160800
rect 82634 159200 82690 160800
rect 82818 159200 82874 160800
rect 83002 159200 83058 160800
rect 83186 159200 83242 160800
rect 83370 159200 83426 160800
rect 83554 159200 83610 160800
rect 83738 159200 83794 160800
rect 83922 159200 83978 160800
rect 84106 159200 84162 160800
rect 84290 159200 84346 160800
rect 84474 159200 84530 160800
rect 84658 159200 84714 160800
rect 84842 159200 84898 160800
rect 110 -800 166 800
rect 294 -800 350 800
rect 478 -800 534 800
rect 662 -800 718 800
rect 846 -800 902 800
rect 1030 -800 1086 800
rect 1214 -800 1270 800
rect 1398 -800 1454 800
rect 1582 -800 1638 800
rect 1766 -800 1822 800
rect 1950 -800 2006 800
rect 2134 -800 2190 800
rect 2318 -800 2374 800
rect 2502 -800 2558 800
rect 2686 -800 2742 800
rect 2870 -800 2926 800
rect 3054 -800 3110 800
rect 3238 -800 3294 800
rect 3422 -800 3478 800
rect 3606 -800 3662 800
rect 3790 -800 3846 800
rect 3974 -800 4030 800
rect 4158 -800 4214 800
rect 4342 -800 4398 800
rect 4526 -800 4582 800
rect 4710 -800 4766 800
rect 4894 -800 4950 800
rect 5078 -800 5134 800
rect 5262 -800 5318 800
rect 5446 -800 5502 800
rect 5630 -800 5686 800
rect 5814 -800 5870 800
rect 5998 -800 6054 800
rect 6182 -800 6238 800
rect 6366 -800 6422 800
rect 6550 -800 6606 800
rect 6734 -800 6790 800
rect 6918 -800 6974 800
rect 7102 -800 7158 800
rect 7286 -800 7342 800
rect 7470 -800 7526 800
rect 7654 -800 7710 800
rect 7838 -800 7894 800
rect 8022 -800 8078 800
rect 8206 -800 8262 800
rect 8390 -800 8446 800
rect 8574 -800 8630 800
rect 8758 -800 8814 800
rect 8942 -800 8998 800
rect 9126 -800 9182 800
rect 9310 -800 9366 800
rect 9494 -800 9550 800
rect 9678 -800 9734 800
rect 9862 -800 9918 800
rect 10046 -800 10102 800
rect 10230 -800 10286 800
rect 10414 -800 10470 800
rect 10598 -800 10654 800
rect 10782 -800 10838 800
rect 10966 -800 11022 800
rect 11150 -800 11206 800
rect 20074 -800 20130 800
rect 20442 -800 20498 800
rect 20810 -800 20866 800
rect 21178 -800 21234 800
rect 21546 -800 21602 800
rect 21914 -800 21970 800
rect 60094 -800 60150 800
rect 60278 -800 60334 800
rect 60462 -800 60518 800
rect 60646 -800 60702 800
rect 60830 -800 60886 800
rect 61014 -800 61070 800
rect 61198 -800 61254 800
rect 61382 -800 61438 800
rect 61566 -800 61622 800
rect 61750 -800 61806 800
rect 61934 -800 61990 800
rect 62118 -800 62174 800
rect 62302 -800 62358 800
rect 62486 -800 62542 800
rect 62670 -800 62726 800
rect 62854 -800 62910 800
rect 63038 -800 63094 800
rect 63222 -800 63278 800
rect 63406 -800 63462 800
rect 63590 -800 63646 800
rect 63774 -800 63830 800
rect 63958 -800 64014 800
rect 64142 -800 64198 800
rect 64326 -800 64382 800
rect 64510 -800 64566 800
rect 64694 -800 64750 800
rect 64878 -800 64934 800
rect 65062 -800 65118 800
rect 65246 -800 65302 800
rect 65430 -800 65486 800
rect 65614 -800 65670 800
rect 65798 -800 65854 800
rect 65982 -800 66038 800
<< obsm2 >>
rect 20 159144 54 159610
rect 222 159144 238 159610
rect 406 159144 422 159610
rect 590 159144 606 159610
rect 774 159144 790 159610
rect 958 159144 974 159610
rect 1142 159144 1158 159610
rect 1326 159144 1342 159610
rect 1510 159144 1526 159610
rect 1694 159144 1710 159610
rect 1878 159144 1894 159610
rect 2062 159144 2078 159610
rect 2246 159144 2262 159610
rect 2430 159144 2446 159610
rect 2614 159144 2630 159610
rect 2798 159144 2814 159610
rect 2982 159144 2998 159610
rect 3166 159144 3182 159610
rect 3350 159144 3366 159610
rect 3534 159144 3550 159610
rect 3718 159144 3734 159610
rect 3902 159144 3918 159610
rect 4086 159144 4102 159610
rect 4270 159144 4286 159610
rect 4454 159144 4470 159610
rect 4638 159144 4654 159610
rect 4822 159144 4838 159610
rect 5006 159144 5022 159610
rect 5190 159144 5206 159610
rect 5374 159144 5390 159610
rect 5558 159144 5574 159610
rect 5742 159144 5758 159610
rect 5926 159144 5942 159610
rect 6110 159144 6126 159610
rect 6294 159144 6310 159610
rect 6478 159144 6494 159610
rect 6662 159144 6678 159610
rect 6846 159144 6862 159610
rect 7030 159144 7046 159610
rect 7214 159144 7230 159610
rect 7398 159144 7414 159610
rect 7582 159144 7598 159610
rect 7766 159144 30046 159610
rect 30214 159144 30230 159610
rect 30398 159144 30414 159610
rect 30582 159144 30598 159610
rect 30766 159144 30782 159610
rect 30950 159144 30966 159610
rect 31134 159144 31150 159610
rect 31318 159144 31334 159610
rect 31502 159144 31518 159610
rect 31686 159144 39982 159610
rect 40150 159144 40166 159610
rect 40334 159144 40350 159610
rect 40518 159144 40534 159610
rect 40702 159144 40718 159610
rect 40886 159144 40902 159610
rect 41070 159144 41086 159610
rect 41254 159144 41270 159610
rect 41438 159144 41454 159610
rect 41622 159144 41638 159610
rect 41806 159144 41822 159610
rect 41990 159144 42006 159610
rect 42174 159144 42190 159610
rect 42358 159144 42374 159610
rect 42542 159144 42558 159610
rect 42726 159144 42742 159610
rect 42910 159144 42926 159610
rect 43094 159144 43110 159610
rect 43278 159144 43294 159610
rect 43462 159144 43478 159610
rect 43646 159144 43662 159610
rect 43830 159144 43846 159610
rect 44014 159144 44030 159610
rect 44198 159144 44214 159610
rect 44382 159144 44398 159610
rect 44566 159144 44582 159610
rect 44750 159144 44766 159610
rect 44934 159144 44950 159610
rect 45118 159144 45134 159610
rect 45302 159144 45318 159610
rect 45486 159144 45502 159610
rect 45670 159144 45686 159610
rect 45854 159144 45870 159610
rect 46038 159144 46054 159610
rect 46222 159144 46238 159610
rect 46406 159144 46422 159610
rect 46590 159144 46606 159610
rect 46774 159144 46790 159610
rect 46958 159144 46974 159610
rect 47142 159144 47158 159610
rect 47326 159144 47342 159610
rect 47510 159144 47526 159610
rect 47694 159144 47710 159610
rect 47878 159144 47894 159610
rect 48062 159144 48078 159610
rect 48246 159144 48262 159610
rect 48430 159144 48446 159610
rect 48614 159144 48630 159610
rect 48798 159144 48814 159610
rect 48982 159144 48998 159610
rect 49166 159144 49182 159610
rect 49350 159144 49366 159610
rect 49534 159144 49550 159610
rect 49718 159144 49734 159610
rect 49902 159144 49918 159610
rect 50086 159144 50102 159610
rect 50270 159144 50286 159610
rect 50454 159144 50470 159610
rect 50638 159144 50654 159610
rect 50822 159144 50838 159610
rect 51006 159144 51022 159610
rect 51190 159144 51206 159610
rect 51374 159144 51390 159610
rect 51558 159144 51574 159610
rect 51742 159144 51758 159610
rect 51926 159144 51942 159610
rect 52110 159144 52126 159610
rect 52294 159144 52310 159610
rect 52478 159144 52494 159610
rect 52662 159144 52678 159610
rect 52846 159144 52862 159610
rect 53030 159144 53046 159610
rect 53214 159144 53230 159610
rect 53398 159144 53414 159610
rect 53582 159144 53598 159610
rect 53766 159144 53782 159610
rect 53950 159144 53966 159610
rect 54134 159144 54150 159610
rect 54318 159144 54334 159610
rect 54502 159144 54518 159610
rect 54686 159144 54702 159610
rect 54870 159144 54886 159610
rect 55054 159144 60038 159610
rect 60206 159144 60222 159610
rect 60390 159144 60406 159610
rect 60574 159144 60590 159610
rect 60758 159144 60774 159610
rect 60942 159144 60958 159610
rect 61126 159144 61142 159610
rect 61310 159144 61326 159610
rect 61494 159144 61510 159610
rect 61678 159144 61694 159610
rect 61862 159144 61878 159610
rect 62046 159144 62062 159610
rect 62230 159144 62246 159610
rect 62414 159144 62430 159610
rect 62598 159144 62614 159610
rect 62782 159144 62798 159610
rect 62966 159144 62982 159610
rect 63150 159144 63166 159610
rect 63334 159144 63350 159610
rect 63518 159144 63534 159610
rect 63702 159144 63718 159610
rect 63886 159144 63902 159610
rect 64070 159144 64086 159610
rect 64254 159144 64270 159610
rect 64438 159144 64454 159610
rect 64622 159144 64638 159610
rect 64806 159144 64822 159610
rect 64990 159144 65006 159610
rect 65174 159144 65190 159610
rect 65358 159144 65374 159610
rect 65542 159144 65558 159610
rect 65726 159144 65742 159610
rect 65910 159144 65926 159610
rect 66094 159144 66110 159610
rect 66278 159144 80002 159610
rect 80170 159144 80186 159610
rect 80354 159144 80370 159610
rect 80538 159144 80554 159610
rect 80722 159144 80738 159610
rect 80906 159144 80922 159610
rect 81090 159144 81106 159610
rect 81274 159144 81290 159610
rect 81458 159144 81474 159610
rect 81642 159144 81658 159610
rect 81826 159144 81842 159610
rect 82010 159144 82026 159610
rect 82194 159144 82210 159610
rect 82378 159144 82394 159610
rect 82562 159144 82578 159610
rect 82746 159144 82762 159610
rect 82930 159144 82946 159610
rect 83114 159144 83130 159610
rect 83298 159144 83314 159610
rect 83482 159144 83498 159610
rect 83666 159144 83682 159610
rect 83850 159144 83866 159610
rect 84034 159144 84050 159610
rect 84218 159144 84234 159610
rect 84402 159144 84418 159610
rect 84586 159144 84602 159610
rect 84770 159144 84786 159610
rect 84954 159144 103114 159610
rect 20 856 103114 159144
rect 20 2 54 856
rect 222 2 238 856
rect 406 2 422 856
rect 590 2 606 856
rect 774 2 790 856
rect 958 2 974 856
rect 1142 2 1158 856
rect 1326 2 1342 856
rect 1510 2 1526 856
rect 1694 2 1710 856
rect 1878 2 1894 856
rect 2062 2 2078 856
rect 2246 2 2262 856
rect 2430 2 2446 856
rect 2614 2 2630 856
rect 2798 2 2814 856
rect 2982 2 2998 856
rect 3166 2 3182 856
rect 3350 2 3366 856
rect 3534 2 3550 856
rect 3718 2 3734 856
rect 3902 2 3918 856
rect 4086 2 4102 856
rect 4270 2 4286 856
rect 4454 2 4470 856
rect 4638 2 4654 856
rect 4822 2 4838 856
rect 5006 2 5022 856
rect 5190 2 5206 856
rect 5374 2 5390 856
rect 5558 2 5574 856
rect 5742 2 5758 856
rect 5926 2 5942 856
rect 6110 2 6126 856
rect 6294 2 6310 856
rect 6478 2 6494 856
rect 6662 2 6678 856
rect 6846 2 6862 856
rect 7030 2 7046 856
rect 7214 2 7230 856
rect 7398 2 7414 856
rect 7582 2 7598 856
rect 7766 2 7782 856
rect 7950 2 7966 856
rect 8134 2 8150 856
rect 8318 2 8334 856
rect 8502 2 8518 856
rect 8686 2 8702 856
rect 8870 2 8886 856
rect 9054 2 9070 856
rect 9238 2 9254 856
rect 9422 2 9438 856
rect 9606 2 9622 856
rect 9790 2 9806 856
rect 9974 2 9990 856
rect 10158 2 10174 856
rect 10342 2 10358 856
rect 10526 2 10542 856
rect 10710 2 10726 856
rect 10894 2 10910 856
rect 11078 2 11094 856
rect 11262 2 20018 856
rect 20186 2 20386 856
rect 20554 2 20754 856
rect 20922 2 21122 856
rect 21290 2 21490 856
rect 21658 2 21858 856
rect 22026 2 60038 856
rect 60206 2 60222 856
rect 60390 2 60406 856
rect 60574 2 60590 856
rect 60758 2 60774 856
rect 60942 2 60958 856
rect 61126 2 61142 856
rect 61310 2 61326 856
rect 61494 2 61510 856
rect 61678 2 61694 856
rect 61862 2 61878 856
rect 62046 2 62062 856
rect 62230 2 62246 856
rect 62414 2 62430 856
rect 62598 2 62614 856
rect 62782 2 62798 856
rect 62966 2 62982 856
rect 63150 2 63166 856
rect 63334 2 63350 856
rect 63518 2 63534 856
rect 63702 2 63718 856
rect 63886 2 63902 856
rect 64070 2 64086 856
rect 64254 2 64270 856
rect 64438 2 64454 856
rect 64622 2 64638 856
rect 64806 2 64822 856
rect 64990 2 65006 856
rect 65174 2 65190 856
rect 65358 2 65374 856
rect 65542 2 65558 856
rect 65726 2 65742 856
rect 65910 2 65926 856
rect 66094 2 103114 856
<< metal3 >>
rect -800 141448 800 141568
rect -800 141176 800 141296
rect -800 140904 800 141024
rect -800 140632 800 140752
rect -800 140360 800 140480
rect -800 140088 800 140208
rect 103200 84056 104800 84176
rect 103200 83512 104800 83632
rect 103200 82968 104800 83088
rect 103200 82424 104800 82544
rect 103200 81880 104800 82000
rect 103200 81336 104800 81456
rect 103200 80792 104800 80912
rect 103200 80248 104800 80368
rect 103200 79704 104800 79824
rect 103200 79160 104800 79280
rect 103200 78616 104800 78736
rect 103200 78072 104800 78192
rect 103200 77528 104800 77648
rect 103200 76984 104800 77104
rect 103200 76440 104800 76560
rect 103200 75896 104800 76016
rect 103200 75352 104800 75472
rect 103200 74808 104800 74928
rect -800 74128 800 74248
rect 103200 74264 104800 74384
rect -800 73856 800 73976
rect -800 73584 800 73704
rect 103200 73720 104800 73840
rect -800 73312 800 73432
rect -800 73040 800 73160
rect 103200 73176 104800 73296
rect -800 72768 800 72888
rect -800 72496 800 72616
rect 103200 72632 104800 72752
rect -800 72224 800 72344
rect -800 71952 800 72072
rect 103200 72088 104800 72208
rect -800 71680 800 71800
rect -800 71408 800 71528
rect 103200 71544 104800 71664
rect -800 71136 800 71256
rect -800 70864 800 70984
rect 103200 71000 104800 71120
rect -800 70592 800 70712
rect -800 70320 800 70440
rect 103200 70456 104800 70576
rect -800 70048 800 70168
rect -800 69776 800 69896
rect 103200 69912 104800 70032
rect -800 69504 800 69624
rect -800 69232 800 69352
rect 103200 69368 104800 69488
rect -800 68960 800 69080
rect -800 68688 800 68808
rect 103200 68824 104800 68944
rect -800 68416 800 68536
rect -800 68144 800 68264
rect 103200 68280 104800 68400
rect -800 67872 800 67992
rect -800 67600 800 67720
rect 103200 67736 104800 67856
rect -800 67328 800 67448
rect -800 67056 800 67176
rect 103200 67192 104800 67312
rect -800 66784 800 66904
rect -800 66512 800 66632
rect 103200 66648 104800 66768
rect -800 66240 800 66360
rect -800 65968 800 66088
rect 103200 66104 104800 66224
rect -800 65696 800 65816
rect -800 65424 800 65544
rect 103200 65560 104800 65680
rect -800 65152 800 65272
rect -800 64880 800 65000
rect 103200 65016 104800 65136
rect -800 64608 800 64728
rect -800 64336 800 64456
rect 103200 64472 104800 64592
rect -800 64064 800 64184
rect -800 63792 800 63912
rect 103200 63928 104800 64048
rect -800 63520 800 63640
rect -800 63248 800 63368
rect 103200 63384 104800 63504
rect -800 62976 800 63096
rect -800 62704 800 62824
rect 103200 62840 104800 62960
rect -800 62432 800 62552
rect -800 62160 800 62280
rect 103200 62296 104800 62416
rect -800 61888 800 62008
rect -800 61616 800 61736
rect 103200 61752 104800 61872
rect -800 61344 800 61464
rect -800 61072 800 61192
rect 103200 61208 104800 61328
rect -800 60800 800 60920
rect -800 60528 800 60648
rect 103200 60664 104800 60784
rect -800 60256 800 60376
rect -800 59984 800 60104
rect 103200 60120 104800 60240
rect -800 59712 800 59832
rect -800 59440 800 59560
rect -800 59168 800 59288
rect -800 58896 800 59016
rect -800 58624 800 58744
rect -800 58352 800 58472
rect -800 58080 800 58200
rect -800 57808 800 57928
rect -800 57536 800 57656
rect -800 57264 800 57384
rect -800 56992 800 57112
rect -800 56720 800 56840
rect -800 56448 800 56568
rect -800 56176 800 56296
rect -800 55904 800 56024
rect -800 55632 800 55752
rect -800 55360 800 55480
rect -800 55088 800 55208
rect -800 54816 800 54936
rect -800 54544 800 54664
rect -800 54272 800 54392
rect -800 54000 800 54120
rect -800 53728 800 53848
rect -800 53456 800 53576
rect -800 53184 800 53304
rect -800 52912 800 53032
rect -800 52640 800 52760
rect -800 52368 800 52488
rect -800 52096 800 52216
rect -800 50736 800 50856
rect -800 50464 800 50584
rect -800 50192 800 50312
rect -800 49920 800 50040
rect -800 49648 800 49768
rect -800 49376 800 49496
rect -800 49104 800 49224
rect -800 48832 800 48952
rect -800 48560 800 48680
rect -800 48288 800 48408
rect -800 48016 800 48136
rect -800 47744 800 47864
rect -800 47472 800 47592
rect -800 47200 800 47320
rect -800 46928 800 47048
rect -800 46656 800 46776
rect -800 46384 800 46504
rect -800 46112 800 46232
rect -800 45840 800 45960
rect -800 45568 800 45688
rect -800 45296 800 45416
rect -800 45024 800 45144
rect -800 44752 800 44872
rect -800 44480 800 44600
rect -800 44208 800 44328
rect -800 43936 800 44056
rect -800 43664 800 43784
rect -800 43392 800 43512
rect -800 43120 800 43240
rect -800 42848 800 42968
rect -800 42576 800 42696
rect -800 42304 800 42424
rect -800 42032 800 42152
rect -800 41760 800 41880
rect -800 41488 800 41608
rect -800 41216 800 41336
rect -800 40944 800 41064
rect -800 40672 800 40792
rect -800 40400 800 40520
rect -800 40128 800 40248
rect -800 18640 800 18760
rect -800 18368 800 18488
rect -800 18096 800 18216
rect -800 17824 800 17944
rect -800 17552 800 17672
rect -800 17280 800 17400
rect -800 17008 800 17128
rect -800 16736 800 16856
rect -800 16464 800 16584
rect -800 16192 800 16312
rect -800 15920 800 16040
rect -800 15648 800 15768
rect -800 15376 800 15496
rect -800 15104 800 15224
rect -800 14832 800 14952
rect -800 14560 800 14680
rect -800 14288 800 14408
rect -800 14016 800 14136
rect -800 13744 800 13864
rect -800 13472 800 13592
rect -800 13200 800 13320
rect -800 12928 800 13048
rect -800 12656 800 12776
rect -800 12384 800 12504
rect -800 12112 800 12232
rect -800 11840 800 11960
rect -800 11568 800 11688
rect -800 11296 800 11416
rect -800 11024 800 11144
rect -800 10752 800 10872
rect -800 10480 800 10600
rect -800 10208 800 10328
rect -800 9936 800 10056
rect -800 9664 800 9784
rect -800 9392 800 9512
rect -800 9120 800 9240
rect -800 8848 800 8968
rect -800 8576 800 8696
rect -800 8304 800 8424
rect -800 8032 800 8152
rect -800 7760 800 7880
rect -800 7488 800 7608
rect -800 7216 800 7336
rect -800 6944 800 7064
rect -800 6672 800 6792
rect -800 6400 800 6520
rect -800 6128 800 6248
rect -800 5856 800 5976
rect -800 5584 800 5704
rect -800 5312 800 5432
rect -800 5040 800 5160
rect -800 4768 800 4888
rect -800 4496 800 4616
rect -800 4224 800 4344
rect -800 3952 800 4072
rect -800 3680 800 3800
rect -800 3408 800 3528
rect -800 3136 800 3256
rect -800 2864 800 2984
rect -800 2592 800 2712
rect -800 2320 800 2440
rect -800 2048 800 2168
rect -800 1776 800 1896
rect -800 1504 800 1624
rect -800 1232 800 1352
rect -800 960 800 1080
rect -800 688 800 808
rect -800 416 800 536
rect -800 144 800 264
rect 103200 4496 104800 4616
rect 103200 4224 104800 4344
rect 103200 3952 104800 4072
rect 103200 3680 104800 3800
rect 103200 3408 104800 3528
rect 103200 3136 104800 3256
rect 103200 2864 104800 2984
rect 103200 2592 104800 2712
rect 103200 2320 104800 2440
rect 103200 2048 104800 2168
rect 103200 1776 104800 1896
rect 103200 1504 104800 1624
rect 103200 1232 104800 1352
rect 103200 960 104800 1080
rect 103200 688 104800 808
rect 103200 416 104800 536
rect 103200 144 104800 264
<< obsm3 >>
rect 197 141648 103200 157793
rect 880 140008 103200 141648
rect 197 84256 103200 140008
rect 197 83976 103120 84256
rect 197 83712 103200 83976
rect 197 83432 103120 83712
rect 197 83168 103200 83432
rect 197 82888 103120 83168
rect 197 82624 103200 82888
rect 197 82344 103120 82624
rect 197 82080 103200 82344
rect 197 81800 103120 82080
rect 197 81536 103200 81800
rect 197 81256 103120 81536
rect 197 80992 103200 81256
rect 197 80712 103120 80992
rect 197 80448 103200 80712
rect 197 80168 103120 80448
rect 197 79904 103200 80168
rect 197 79624 103120 79904
rect 197 79360 103200 79624
rect 197 79080 103120 79360
rect 197 78816 103200 79080
rect 197 78536 103120 78816
rect 197 78272 103200 78536
rect 197 77992 103120 78272
rect 197 77728 103200 77992
rect 197 77448 103120 77728
rect 197 77184 103200 77448
rect 197 76904 103120 77184
rect 197 76640 103200 76904
rect 197 76360 103120 76640
rect 197 76096 103200 76360
rect 197 75816 103120 76096
rect 197 75552 103200 75816
rect 197 75272 103120 75552
rect 197 75008 103200 75272
rect 197 74728 103120 75008
rect 197 74464 103200 74728
rect 197 74328 103120 74464
rect 880 74184 103120 74328
rect 880 73920 103200 74184
rect 880 73640 103120 73920
rect 880 73376 103200 73640
rect 880 73096 103120 73376
rect 880 72832 103200 73096
rect 880 72552 103120 72832
rect 880 72288 103200 72552
rect 880 72008 103120 72288
rect 880 71744 103200 72008
rect 880 71464 103120 71744
rect 880 71200 103200 71464
rect 880 70920 103120 71200
rect 880 70656 103200 70920
rect 880 70376 103120 70656
rect 880 70112 103200 70376
rect 880 69832 103120 70112
rect 880 69568 103200 69832
rect 880 69288 103120 69568
rect 880 69024 103200 69288
rect 880 68744 103120 69024
rect 880 68480 103200 68744
rect 880 68200 103120 68480
rect 880 67936 103200 68200
rect 880 67656 103120 67936
rect 880 67392 103200 67656
rect 880 67112 103120 67392
rect 880 66848 103200 67112
rect 880 66568 103120 66848
rect 880 66304 103200 66568
rect 880 66024 103120 66304
rect 880 65760 103200 66024
rect 880 65480 103120 65760
rect 880 65216 103200 65480
rect 880 64936 103120 65216
rect 880 64672 103200 64936
rect 880 64392 103120 64672
rect 880 64128 103200 64392
rect 880 63848 103120 64128
rect 880 63584 103200 63848
rect 880 63304 103120 63584
rect 880 63040 103200 63304
rect 880 62760 103120 63040
rect 880 62496 103200 62760
rect 880 62216 103120 62496
rect 880 61952 103200 62216
rect 880 61672 103120 61952
rect 880 61408 103200 61672
rect 880 61128 103120 61408
rect 880 60864 103200 61128
rect 880 60584 103120 60864
rect 880 60320 103200 60584
rect 880 60040 103120 60320
rect 880 52016 103200 60040
rect 197 50936 103200 52016
rect 880 40048 103200 50936
rect 197 18840 103200 40048
rect 880 4696 103200 18840
rect 880 171 103120 4696
<< metal4 >>
rect 3748 2128 4988 157808
rect 13748 2128 14988 157808
rect 23748 2128 24988 157808
rect 33748 2128 34988 157808
rect 43748 2128 44988 157808
rect 53748 2128 54988 157808
rect 63748 2128 64988 157808
rect 73748 2128 74988 157808
rect 83748 2128 84988 157808
rect 93748 2128 94988 157808
<< obsm4 >>
rect 243 2048 3668 157589
rect 5068 2048 13668 157589
rect 15068 2048 23668 157589
rect 25068 2048 33668 157589
rect 35068 2048 43668 157589
rect 45068 2048 53668 157589
rect 55068 2048 63668 157589
rect 65068 2048 73668 157589
rect 75068 2048 83668 157589
rect 85068 2048 89733 157589
rect 243 715 89733 2048
<< labels >>
rlabel metal3 s -800 49920 800 50040 4 cfg_cska_pinmux[0]
port 1 nsew signal input
rlabel metal3 s -800 49648 800 49768 4 cfg_cska_pinmux[1]
port 2 nsew signal input
rlabel metal3 s -800 49376 800 49496 4 cfg_cska_pinmux[2]
port 3 nsew signal input
rlabel metal3 s -800 49104 800 49224 4 cfg_cska_pinmux[3]
port 4 nsew signal input
rlabel metal2 s 66166 159200 66222 160800 6 cfg_dc_trim[0]
port 5 nsew signal output
rlabel metal2 s 64326 159200 64382 160800 6 cfg_dc_trim[10]
port 6 nsew signal output
rlabel metal2 s 64142 159200 64198 160800 6 cfg_dc_trim[11]
port 7 nsew signal output
rlabel metal2 s 63958 159200 64014 160800 6 cfg_dc_trim[12]
port 8 nsew signal output
rlabel metal2 s 63774 159200 63830 160800 6 cfg_dc_trim[13]
port 9 nsew signal output
rlabel metal2 s 63590 159200 63646 160800 6 cfg_dc_trim[14]
port 10 nsew signal output
rlabel metal2 s 63406 159200 63462 160800 6 cfg_dc_trim[15]
port 11 nsew signal output
rlabel metal2 s 63222 159200 63278 160800 6 cfg_dc_trim[16]
port 12 nsew signal output
rlabel metal2 s 63038 159200 63094 160800 6 cfg_dc_trim[17]
port 13 nsew signal output
rlabel metal2 s 62854 159200 62910 160800 6 cfg_dc_trim[18]
port 14 nsew signal output
rlabel metal2 s 62670 159200 62726 160800 6 cfg_dc_trim[19]
port 15 nsew signal output
rlabel metal2 s 65982 159200 66038 160800 6 cfg_dc_trim[1]
port 16 nsew signal output
rlabel metal2 s 62486 159200 62542 160800 6 cfg_dc_trim[20]
port 17 nsew signal output
rlabel metal2 s 62302 159200 62358 160800 6 cfg_dc_trim[21]
port 18 nsew signal output
rlabel metal2 s 62118 159200 62174 160800 6 cfg_dc_trim[22]
port 19 nsew signal output
rlabel metal2 s 61934 159200 61990 160800 6 cfg_dc_trim[23]
port 20 nsew signal output
rlabel metal2 s 61750 159200 61806 160800 6 cfg_dc_trim[24]
port 21 nsew signal output
rlabel metal2 s 61566 159200 61622 160800 6 cfg_dc_trim[25]
port 22 nsew signal output
rlabel metal2 s 65798 159200 65854 160800 6 cfg_dc_trim[2]
port 23 nsew signal output
rlabel metal2 s 65614 159200 65670 160800 6 cfg_dc_trim[3]
port 24 nsew signal output
rlabel metal2 s 65430 159200 65486 160800 6 cfg_dc_trim[4]
port 25 nsew signal output
rlabel metal2 s 65246 159200 65302 160800 6 cfg_dc_trim[5]
port 26 nsew signal output
rlabel metal2 s 65062 159200 65118 160800 6 cfg_dc_trim[6]
port 27 nsew signal output
rlabel metal2 s 64878 159200 64934 160800 6 cfg_dc_trim[7]
port 28 nsew signal output
rlabel metal2 s 64694 159200 64750 160800 6 cfg_dc_trim[8]
port 29 nsew signal output
rlabel metal2 s 64510 159200 64566 160800 6 cfg_dc_trim[9]
port 30 nsew signal output
rlabel metal2 s 60094 159200 60150 160800 6 cfg_dco_mode
port 31 nsew signal output
rlabel metal2 s 60278 159200 60334 160800 6 cfg_pll_enb
port 32 nsew signal output
rlabel metal2 s 61382 159200 61438 160800 6 cfg_pll_fed_div[0]
port 33 nsew signal output
rlabel metal2 s 61198 159200 61254 160800 6 cfg_pll_fed_div[1]
port 34 nsew signal output
rlabel metal2 s 61014 159200 61070 160800 6 cfg_pll_fed_div[2]
port 35 nsew signal output
rlabel metal2 s 60830 159200 60886 160800 6 cfg_pll_fed_div[3]
port 36 nsew signal output
rlabel metal2 s 60646 159200 60702 160800 6 cfg_pll_fed_div[4]
port 37 nsew signal output
rlabel metal2 s 4894 -800 4950 800 8 cfg_riscv_ctrl[0]
port 38 nsew signal output
rlabel metal2 s 3054 -800 3110 800 8 cfg_riscv_ctrl[10]
port 39 nsew signal output
rlabel metal2 s 2870 -800 2926 800 8 cfg_riscv_ctrl[11]
port 40 nsew signal output
rlabel metal2 s 2686 -800 2742 800 8 cfg_riscv_ctrl[12]
port 41 nsew signal output
rlabel metal2 s 2502 -800 2558 800 8 cfg_riscv_ctrl[13]
port 42 nsew signal output
rlabel metal2 s 2318 -800 2374 800 8 cfg_riscv_ctrl[14]
port 43 nsew signal output
rlabel metal2 s 2134 -800 2190 800 8 cfg_riscv_ctrl[15]
port 44 nsew signal output
rlabel metal2 s 4710 -800 4766 800 8 cfg_riscv_ctrl[1]
port 45 nsew signal output
rlabel metal2 s 4526 -800 4582 800 8 cfg_riscv_ctrl[2]
port 46 nsew signal output
rlabel metal2 s 4342 -800 4398 800 8 cfg_riscv_ctrl[3]
port 47 nsew signal output
rlabel metal2 s 4158 -800 4214 800 8 cfg_riscv_ctrl[4]
port 48 nsew signal output
rlabel metal2 s 3974 -800 4030 800 8 cfg_riscv_ctrl[5]
port 49 nsew signal output
rlabel metal2 s 3790 -800 3846 800 8 cfg_riscv_ctrl[6]
port 50 nsew signal output
rlabel metal2 s 3606 -800 3662 800 8 cfg_riscv_ctrl[7]
port 51 nsew signal output
rlabel metal2 s 3422 -800 3478 800 8 cfg_riscv_ctrl[8]
port 52 nsew signal output
rlabel metal2 s 3238 -800 3294 800 8 cfg_riscv_ctrl[9]
port 53 nsew signal output
rlabel metal3 s -800 18640 800 18760 4 cfg_strap_pad_ctrl
port 54 nsew signal input
rlabel metal2 s 65982 -800 66038 800 8 cpu_clk
port 55 nsew signal input
rlabel metal2 s 662 -800 718 800 8 cpu_core_rst_n[0]
port 56 nsew signal output
rlabel metal2 s 478 -800 534 800 8 cpu_core_rst_n[1]
port 57 nsew signal output
rlabel metal2 s 294 -800 350 800 8 cpu_core_rst_n[2]
port 58 nsew signal output
rlabel metal2 s 110 -800 166 800 8 cpu_core_rst_n[3]
port 59 nsew signal output
rlabel metal2 s 846 -800 902 800 8 cpu_intf_rst_n
port 60 nsew signal output
rlabel metal3 s 103200 60120 104800 60240 6 digital_io_in[0]
port 61 nsew signal input
rlabel metal3 s 103200 76440 104800 76560 6 digital_io_in[10]
port 62 nsew signal input
rlabel metal3 s 103200 78072 104800 78192 6 digital_io_in[11]
port 63 nsew signal input
rlabel metal3 s 103200 79704 104800 79824 6 digital_io_in[12]
port 64 nsew signal input
rlabel metal3 s 103200 81336 104800 81456 6 digital_io_in[13]
port 65 nsew signal input
rlabel metal3 s 103200 82968 104800 83088 6 digital_io_in[14]
port 66 nsew signal input
rlabel metal2 s 84474 159200 84530 160800 6 digital_io_in[15]
port 67 nsew signal input
rlabel metal2 s 83922 159200 83978 160800 6 digital_io_in[16]
port 68 nsew signal input
rlabel metal2 s 83370 159200 83426 160800 6 digital_io_in[17]
port 69 nsew signal input
rlabel metal2 s 82818 159200 82874 160800 6 digital_io_in[18]
port 70 nsew signal input
rlabel metal2 s 82266 159200 82322 160800 6 digital_io_in[19]
port 71 nsew signal input
rlabel metal3 s 103200 61752 104800 61872 6 digital_io_in[1]
port 72 nsew signal input
rlabel metal2 s 81714 159200 81770 160800 6 digital_io_in[20]
port 73 nsew signal input
rlabel metal2 s 81162 159200 81218 160800 6 digital_io_in[21]
port 74 nsew signal input
rlabel metal2 s 80610 159200 80666 160800 6 digital_io_in[22]
port 75 nsew signal input
rlabel metal2 s 80058 159200 80114 160800 6 digital_io_in[23]
port 76 nsew signal input
rlabel metal2 s 7654 159200 7710 160800 6 digital_io_in[24]
port 77 nsew signal input
rlabel metal2 s 7102 159200 7158 160800 6 digital_io_in[25]
port 78 nsew signal input
rlabel metal2 s 6550 159200 6606 160800 6 digital_io_in[26]
port 79 nsew signal input
rlabel metal2 s 5998 159200 6054 160800 6 digital_io_in[27]
port 80 nsew signal input
rlabel metal2 s 5446 159200 5502 160800 6 digital_io_in[28]
port 81 nsew signal input
rlabel metal2 s 4894 159200 4950 160800 6 digital_io_in[29]
port 82 nsew signal input
rlabel metal3 s 103200 63384 104800 63504 6 digital_io_in[2]
port 83 nsew signal input
rlabel metal2 s 4342 159200 4398 160800 6 digital_io_in[30]
port 84 nsew signal input
rlabel metal2 s 3790 159200 3846 160800 6 digital_io_in[31]
port 85 nsew signal input
rlabel metal2 s 3238 159200 3294 160800 6 digital_io_in[32]
port 86 nsew signal input
rlabel metal2 s 2686 159200 2742 160800 6 digital_io_in[33]
port 87 nsew signal input
rlabel metal2 s 2134 159200 2190 160800 6 digital_io_in[34]
port 88 nsew signal input
rlabel metal2 s 1582 159200 1638 160800 6 digital_io_in[35]
port 89 nsew signal input
rlabel metal2 s 1030 159200 1086 160800 6 digital_io_in[36]
port 90 nsew signal input
rlabel metal2 s 478 159200 534 160800 6 digital_io_in[37]
port 91 nsew signal input
rlabel metal3 s 103200 65016 104800 65136 6 digital_io_in[3]
port 92 nsew signal input
rlabel metal3 s 103200 66648 104800 66768 6 digital_io_in[4]
port 93 nsew signal input
rlabel metal3 s 103200 68280 104800 68400 6 digital_io_in[5]
port 94 nsew signal input
rlabel metal3 s 103200 69912 104800 70032 6 digital_io_in[6]
port 95 nsew signal input
rlabel metal3 s 103200 71544 104800 71664 6 digital_io_in[7]
port 96 nsew signal input
rlabel metal3 s 103200 73176 104800 73296 6 digital_io_in[8]
port 97 nsew signal input
rlabel metal3 s 103200 74808 104800 74928 6 digital_io_in[9]
port 98 nsew signal input
rlabel metal3 s 103200 61208 104800 61328 6 digital_io_oen[0]
port 99 nsew signal output
rlabel metal3 s 103200 77528 104800 77648 6 digital_io_oen[10]
port 100 nsew signal output
rlabel metal3 s 103200 79160 104800 79280 6 digital_io_oen[11]
port 101 nsew signal output
rlabel metal3 s 103200 80792 104800 80912 6 digital_io_oen[12]
port 102 nsew signal output
rlabel metal3 s 103200 82424 104800 82544 6 digital_io_oen[13]
port 103 nsew signal output
rlabel metal3 s 103200 84056 104800 84176 6 digital_io_oen[14]
port 104 nsew signal output
rlabel metal2 s 84842 159200 84898 160800 6 digital_io_oen[15]
port 105 nsew signal output
rlabel metal2 s 84290 159200 84346 160800 6 digital_io_oen[16]
port 106 nsew signal output
rlabel metal2 s 83738 159200 83794 160800 6 digital_io_oen[17]
port 107 nsew signal output
rlabel metal2 s 83186 159200 83242 160800 6 digital_io_oen[18]
port 108 nsew signal output
rlabel metal2 s 82634 159200 82690 160800 6 digital_io_oen[19]
port 109 nsew signal output
rlabel metal3 s 103200 62840 104800 62960 6 digital_io_oen[1]
port 110 nsew signal output
rlabel metal2 s 82082 159200 82138 160800 6 digital_io_oen[20]
port 111 nsew signal output
rlabel metal2 s 81530 159200 81586 160800 6 digital_io_oen[21]
port 112 nsew signal output
rlabel metal2 s 80978 159200 81034 160800 6 digital_io_oen[22]
port 113 nsew signal output
rlabel metal2 s 80426 159200 80482 160800 6 digital_io_oen[23]
port 114 nsew signal output
rlabel metal2 s 7286 159200 7342 160800 6 digital_io_oen[24]
port 115 nsew signal output
rlabel metal2 s 6734 159200 6790 160800 6 digital_io_oen[25]
port 116 nsew signal output
rlabel metal2 s 6182 159200 6238 160800 6 digital_io_oen[26]
port 117 nsew signal output
rlabel metal2 s 5630 159200 5686 160800 6 digital_io_oen[27]
port 118 nsew signal output
rlabel metal2 s 5078 159200 5134 160800 6 digital_io_oen[28]
port 119 nsew signal output
rlabel metal2 s 4526 159200 4582 160800 6 digital_io_oen[29]
port 120 nsew signal output
rlabel metal3 s 103200 64472 104800 64592 6 digital_io_oen[2]
port 121 nsew signal output
rlabel metal2 s 3974 159200 4030 160800 6 digital_io_oen[30]
port 122 nsew signal output
rlabel metal2 s 3422 159200 3478 160800 6 digital_io_oen[31]
port 123 nsew signal output
rlabel metal2 s 2870 159200 2926 160800 6 digital_io_oen[32]
port 124 nsew signal output
rlabel metal2 s 2318 159200 2374 160800 6 digital_io_oen[33]
port 125 nsew signal output
rlabel metal2 s 1766 159200 1822 160800 6 digital_io_oen[34]
port 126 nsew signal output
rlabel metal2 s 1214 159200 1270 160800 6 digital_io_oen[35]
port 127 nsew signal output
rlabel metal2 s 662 159200 718 160800 6 digital_io_oen[36]
port 128 nsew signal output
rlabel metal2 s 110 159200 166 160800 6 digital_io_oen[37]
port 129 nsew signal output
rlabel metal3 s 103200 66104 104800 66224 6 digital_io_oen[3]
port 130 nsew signal output
rlabel metal3 s 103200 67736 104800 67856 6 digital_io_oen[4]
port 131 nsew signal output
rlabel metal3 s 103200 69368 104800 69488 6 digital_io_oen[5]
port 132 nsew signal output
rlabel metal3 s 103200 71000 104800 71120 6 digital_io_oen[6]
port 133 nsew signal output
rlabel metal3 s 103200 72632 104800 72752 6 digital_io_oen[7]
port 134 nsew signal output
rlabel metal3 s 103200 74264 104800 74384 6 digital_io_oen[8]
port 135 nsew signal output
rlabel metal3 s 103200 75896 104800 76016 6 digital_io_oen[9]
port 136 nsew signal output
rlabel metal3 s 103200 60664 104800 60784 6 digital_io_out[0]
port 137 nsew signal output
rlabel metal3 s 103200 76984 104800 77104 6 digital_io_out[10]
port 138 nsew signal output
rlabel metal3 s 103200 78616 104800 78736 6 digital_io_out[11]
port 139 nsew signal output
rlabel metal3 s 103200 80248 104800 80368 6 digital_io_out[12]
port 140 nsew signal output
rlabel metal3 s 103200 81880 104800 82000 6 digital_io_out[13]
port 141 nsew signal output
rlabel metal3 s 103200 83512 104800 83632 6 digital_io_out[14]
port 142 nsew signal output
rlabel metal2 s 84658 159200 84714 160800 6 digital_io_out[15]
port 143 nsew signal output
rlabel metal2 s 84106 159200 84162 160800 6 digital_io_out[16]
port 144 nsew signal output
rlabel metal2 s 83554 159200 83610 160800 6 digital_io_out[17]
port 145 nsew signal output
rlabel metal2 s 83002 159200 83058 160800 6 digital_io_out[18]
port 146 nsew signal output
rlabel metal2 s 82450 159200 82506 160800 6 digital_io_out[19]
port 147 nsew signal output
rlabel metal3 s 103200 62296 104800 62416 6 digital_io_out[1]
port 148 nsew signal output
rlabel metal2 s 81898 159200 81954 160800 6 digital_io_out[20]
port 149 nsew signal output
rlabel metal2 s 81346 159200 81402 160800 6 digital_io_out[21]
port 150 nsew signal output
rlabel metal2 s 80794 159200 80850 160800 6 digital_io_out[22]
port 151 nsew signal output
rlabel metal2 s 80242 159200 80298 160800 6 digital_io_out[23]
port 152 nsew signal output
rlabel metal2 s 7470 159200 7526 160800 6 digital_io_out[24]
port 153 nsew signal output
rlabel metal2 s 6918 159200 6974 160800 6 digital_io_out[25]
port 154 nsew signal output
rlabel metal2 s 6366 159200 6422 160800 6 digital_io_out[26]
port 155 nsew signal output
rlabel metal2 s 5814 159200 5870 160800 6 digital_io_out[27]
port 156 nsew signal output
rlabel metal2 s 5262 159200 5318 160800 6 digital_io_out[28]
port 157 nsew signal output
rlabel metal2 s 4710 159200 4766 160800 6 digital_io_out[29]
port 158 nsew signal output
rlabel metal3 s 103200 63928 104800 64048 6 digital_io_out[2]
port 159 nsew signal output
rlabel metal2 s 4158 159200 4214 160800 6 digital_io_out[30]
port 160 nsew signal output
rlabel metal2 s 3606 159200 3662 160800 6 digital_io_out[31]
port 161 nsew signal output
rlabel metal2 s 3054 159200 3110 160800 6 digital_io_out[32]
port 162 nsew signal output
rlabel metal2 s 2502 159200 2558 160800 6 digital_io_out[33]
port 163 nsew signal output
rlabel metal2 s 1950 159200 2006 160800 6 digital_io_out[34]
port 164 nsew signal output
rlabel metal2 s 1398 159200 1454 160800 6 digital_io_out[35]
port 165 nsew signal output
rlabel metal2 s 846 159200 902 160800 6 digital_io_out[36]
port 166 nsew signal output
rlabel metal2 s 294 159200 350 160800 6 digital_io_out[37]
port 167 nsew signal output
rlabel metal3 s 103200 65560 104800 65680 6 digital_io_out[3]
port 168 nsew signal output
rlabel metal3 s 103200 67192 104800 67312 6 digital_io_out[4]
port 169 nsew signal output
rlabel metal3 s 103200 68824 104800 68944 6 digital_io_out[5]
port 170 nsew signal output
rlabel metal3 s 103200 70456 104800 70576 6 digital_io_out[6]
port 171 nsew signal output
rlabel metal3 s 103200 72088 104800 72208 6 digital_io_out[7]
port 172 nsew signal output
rlabel metal3 s 103200 73720 104800 73840 6 digital_io_out[8]
port 173 nsew signal output
rlabel metal3 s 103200 75352 104800 75472 6 digital_io_out[9]
port 174 nsew signal output
rlabel metal3 s -800 18368 800 18488 4 e_reset_n
port 175 nsew signal input
rlabel metal2 s 7470 -800 7526 800 8 i2cm_clk_i
port 176 nsew signal output
rlabel metal2 s 7286 -800 7342 800 8 i2cm_clk_o
port 177 nsew signal input
rlabel metal2 s 7654 -800 7710 800 8 i2cm_clk_oen
port 178 nsew signal input
rlabel metal2 s 8206 -800 8262 800 8 i2cm_data_i
port 179 nsew signal output
rlabel metal2 s 8022 -800 8078 800 8 i2cm_data_o
port 180 nsew signal input
rlabel metal2 s 7838 -800 7894 800 8 i2cm_data_oen
port 181 nsew signal input
rlabel metal2 s 9862 -800 9918 800 8 i2cm_intr
port 182 nsew signal input
rlabel metal2 s 1766 -800 1822 800 8 i2cm_rst_n
port 183 nsew signal output
rlabel metal2 s 20810 -800 20866 800 8 int_pll_clock
port 184 nsew signal input
rlabel metal2 s 30838 159200 30894 160800 6 ir_intr
port 185 nsew signal input
rlabel metal2 s 30470 159200 30526 160800 6 ir_rx
port 186 nsew signal output
rlabel metal2 s 30654 159200 30710 160800 6 ir_tx
port 187 nsew signal input
rlabel metal3 s -800 48832 800 48952 4 irq_lines[0]
port 188 nsew signal output
rlabel metal3 s -800 46112 800 46232 4 irq_lines[10]
port 189 nsew signal output
rlabel metal3 s -800 45840 800 45960 4 irq_lines[11]
port 190 nsew signal output
rlabel metal3 s -800 45568 800 45688 4 irq_lines[12]
port 191 nsew signal output
rlabel metal3 s -800 45296 800 45416 4 irq_lines[13]
port 192 nsew signal output
rlabel metal3 s -800 45024 800 45144 4 irq_lines[14]
port 193 nsew signal output
rlabel metal3 s -800 44752 800 44872 4 irq_lines[15]
port 194 nsew signal output
rlabel metal3 s -800 44480 800 44600 4 irq_lines[16]
port 195 nsew signal output
rlabel metal3 s -800 44208 800 44328 4 irq_lines[17]
port 196 nsew signal output
rlabel metal3 s -800 43936 800 44056 4 irq_lines[18]
port 197 nsew signal output
rlabel metal3 s -800 43664 800 43784 4 irq_lines[19]
port 198 nsew signal output
rlabel metal3 s -800 48560 800 48680 4 irq_lines[1]
port 199 nsew signal output
rlabel metal3 s -800 43392 800 43512 4 irq_lines[20]
port 200 nsew signal output
rlabel metal3 s -800 43120 800 43240 4 irq_lines[21]
port 201 nsew signal output
rlabel metal3 s -800 42848 800 42968 4 irq_lines[22]
port 202 nsew signal output
rlabel metal3 s -800 42576 800 42696 4 irq_lines[23]
port 203 nsew signal output
rlabel metal3 s -800 42304 800 42424 4 irq_lines[24]
port 204 nsew signal output
rlabel metal3 s -800 42032 800 42152 4 irq_lines[25]
port 205 nsew signal output
rlabel metal3 s -800 41760 800 41880 4 irq_lines[26]
port 206 nsew signal output
rlabel metal3 s -800 41488 800 41608 4 irq_lines[27]
port 207 nsew signal output
rlabel metal3 s -800 41216 800 41336 4 irq_lines[28]
port 208 nsew signal output
rlabel metal3 s -800 40944 800 41064 4 irq_lines[29]
port 209 nsew signal output
rlabel metal3 s -800 48288 800 48408 4 irq_lines[2]
port 210 nsew signal output
rlabel metal3 s -800 40672 800 40792 4 irq_lines[30]
port 211 nsew signal output
rlabel metal3 s -800 40400 800 40520 4 irq_lines[31]
port 212 nsew signal output
rlabel metal3 s -800 48016 800 48136 4 irq_lines[3]
port 213 nsew signal output
rlabel metal3 s -800 47744 800 47864 4 irq_lines[4]
port 214 nsew signal output
rlabel metal3 s -800 47472 800 47592 4 irq_lines[5]
port 215 nsew signal output
rlabel metal3 s -800 47200 800 47320 4 irq_lines[6]
port 216 nsew signal output
rlabel metal3 s -800 46928 800 47048 4 irq_lines[7]
port 217 nsew signal output
rlabel metal3 s -800 46656 800 46776 4 irq_lines[8]
port 218 nsew signal output
rlabel metal3 s -800 46384 800 46504 4 irq_lines[9]
port 219 nsew signal output
rlabel metal3 s -800 50736 800 50856 4 mclk
port 220 nsew signal input
rlabel metal3 s -800 18096 800 18216 4 p_reset_n
port 221 nsew signal input
rlabel metal2 s 60094 -800 60150 800 8 pinmux_debug[0]
port 222 nsew signal output
rlabel metal2 s 61934 -800 61990 800 8 pinmux_debug[10]
port 223 nsew signal output
rlabel metal2 s 62118 -800 62174 800 8 pinmux_debug[11]
port 224 nsew signal output
rlabel metal2 s 62302 -800 62358 800 8 pinmux_debug[12]
port 225 nsew signal output
rlabel metal2 s 62486 -800 62542 800 8 pinmux_debug[13]
port 226 nsew signal output
rlabel metal2 s 62670 -800 62726 800 8 pinmux_debug[14]
port 227 nsew signal output
rlabel metal2 s 62854 -800 62910 800 8 pinmux_debug[15]
port 228 nsew signal output
rlabel metal2 s 63038 -800 63094 800 8 pinmux_debug[16]
port 229 nsew signal output
rlabel metal2 s 63222 -800 63278 800 8 pinmux_debug[17]
port 230 nsew signal output
rlabel metal2 s 63406 -800 63462 800 8 pinmux_debug[18]
port 231 nsew signal output
rlabel metal2 s 63590 -800 63646 800 8 pinmux_debug[19]
port 232 nsew signal output
rlabel metal2 s 60278 -800 60334 800 8 pinmux_debug[1]
port 233 nsew signal output
rlabel metal2 s 63774 -800 63830 800 8 pinmux_debug[20]
port 234 nsew signal output
rlabel metal2 s 63958 -800 64014 800 8 pinmux_debug[21]
port 235 nsew signal output
rlabel metal2 s 64142 -800 64198 800 8 pinmux_debug[22]
port 236 nsew signal output
rlabel metal2 s 64326 -800 64382 800 8 pinmux_debug[23]
port 237 nsew signal output
rlabel metal2 s 64510 -800 64566 800 8 pinmux_debug[24]
port 238 nsew signal output
rlabel metal2 s 64694 -800 64750 800 8 pinmux_debug[25]
port 239 nsew signal output
rlabel metal2 s 64878 -800 64934 800 8 pinmux_debug[26]
port 240 nsew signal output
rlabel metal2 s 65062 -800 65118 800 8 pinmux_debug[27]
port 241 nsew signal output
rlabel metal2 s 65246 -800 65302 800 8 pinmux_debug[28]
port 242 nsew signal output
rlabel metal2 s 65430 -800 65486 800 8 pinmux_debug[29]
port 243 nsew signal output
rlabel metal2 s 60462 -800 60518 800 8 pinmux_debug[2]
port 244 nsew signal output
rlabel metal2 s 65614 -800 65670 800 8 pinmux_debug[30]
port 245 nsew signal output
rlabel metal2 s 65798 -800 65854 800 8 pinmux_debug[31]
port 246 nsew signal output
rlabel metal2 s 60646 -800 60702 800 8 pinmux_debug[3]
port 247 nsew signal output
rlabel metal2 s 60830 -800 60886 800 8 pinmux_debug[4]
port 248 nsew signal output
rlabel metal2 s 61014 -800 61070 800 8 pinmux_debug[5]
port 249 nsew signal output
rlabel metal2 s 61198 -800 61254 800 8 pinmux_debug[6]
port 250 nsew signal output
rlabel metal2 s 61382 -800 61438 800 8 pinmux_debug[7]
port 251 nsew signal output
rlabel metal2 s 61566 -800 61622 800 8 pinmux_debug[8]
port 252 nsew signal output
rlabel metal2 s 61750 -800 61806 800 8 pinmux_debug[9]
port 253 nsew signal output
rlabel metal2 s 60462 159200 60518 160800 6 pll_ref_clk
port 254 nsew signal output
rlabel metal2 s 9678 -800 9734 800 8 pulse1m_mclk
port 255 nsew signal output
rlabel metal2 s 1030 -800 1086 800 8 qspim_rst_n
port 256 nsew signal output
rlabel metal3 s -800 74128 800 74248 4 reg_ack
port 257 nsew signal output
rlabel metal3 s -800 55360 800 55480 4 reg_addr[0]
port 258 nsew signal input
rlabel metal3 s -800 52640 800 52760 4 reg_addr[10]
port 259 nsew signal input
rlabel metal3 s -800 55088 800 55208 4 reg_addr[1]
port 260 nsew signal input
rlabel metal3 s -800 54816 800 54936 4 reg_addr[2]
port 261 nsew signal input
rlabel metal3 s -800 54544 800 54664 4 reg_addr[3]
port 262 nsew signal input
rlabel metal3 s -800 54272 800 54392 4 reg_addr[4]
port 263 nsew signal input
rlabel metal3 s -800 54000 800 54120 4 reg_addr[5]
port 264 nsew signal input
rlabel metal3 s -800 53728 800 53848 4 reg_addr[6]
port 265 nsew signal input
rlabel metal3 s -800 53456 800 53576 4 reg_addr[7]
port 266 nsew signal input
rlabel metal3 s -800 53184 800 53304 4 reg_addr[8]
port 267 nsew signal input
rlabel metal3 s -800 52912 800 53032 4 reg_addr[9]
port 268 nsew signal input
rlabel metal3 s -800 56448 800 56568 4 reg_be[0]
port 269 nsew signal input
rlabel metal3 s -800 56176 800 56296 4 reg_be[1]
port 270 nsew signal input
rlabel metal3 s -800 55904 800 56024 4 reg_be[2]
port 271 nsew signal input
rlabel metal3 s -800 55632 800 55752 4 reg_be[3]
port 272 nsew signal input
rlabel metal3 s -800 52096 800 52216 4 reg_cs
port 273 nsew signal input
rlabel metal2 s 54942 159200 54998 160800 6 reg_peri_ack
port 274 nsew signal input
rlabel metal2 s 42246 159200 42302 160800 6 reg_peri_addr[0]
port 275 nsew signal output
rlabel metal2 s 40406 159200 40462 160800 6 reg_peri_addr[10]
port 276 nsew signal output
rlabel metal2 s 42062 159200 42118 160800 6 reg_peri_addr[1]
port 277 nsew signal output
rlabel metal2 s 41878 159200 41934 160800 6 reg_peri_addr[2]
port 278 nsew signal output
rlabel metal2 s 41694 159200 41750 160800 6 reg_peri_addr[3]
port 279 nsew signal output
rlabel metal2 s 41510 159200 41566 160800 6 reg_peri_addr[4]
port 280 nsew signal output
rlabel metal2 s 41326 159200 41382 160800 6 reg_peri_addr[5]
port 281 nsew signal output
rlabel metal2 s 41142 159200 41198 160800 6 reg_peri_addr[6]
port 282 nsew signal output
rlabel metal2 s 40958 159200 41014 160800 6 reg_peri_addr[7]
port 283 nsew signal output
rlabel metal2 s 40774 159200 40830 160800 6 reg_peri_addr[8]
port 284 nsew signal output
rlabel metal2 s 40590 159200 40646 160800 6 reg_peri_addr[9]
port 285 nsew signal output
rlabel metal2 s 42982 159200 43038 160800 6 reg_peri_be[0]
port 286 nsew signal output
rlabel metal2 s 42798 159200 42854 160800 6 reg_peri_be[1]
port 287 nsew signal output
rlabel metal2 s 42614 159200 42670 160800 6 reg_peri_be[2]
port 288 nsew signal output
rlabel metal2 s 42430 159200 42486 160800 6 reg_peri_be[3]
port 289 nsew signal output
rlabel metal2 s 40038 159200 40094 160800 6 reg_peri_cs
port 290 nsew signal output
rlabel metal2 s 54758 159200 54814 160800 6 reg_peri_rdata[0]
port 291 nsew signal input
rlabel metal2 s 52918 159200 52974 160800 6 reg_peri_rdata[10]
port 292 nsew signal input
rlabel metal2 s 52734 159200 52790 160800 6 reg_peri_rdata[11]
port 293 nsew signal input
rlabel metal2 s 52550 159200 52606 160800 6 reg_peri_rdata[12]
port 294 nsew signal input
rlabel metal2 s 52366 159200 52422 160800 6 reg_peri_rdata[13]
port 295 nsew signal input
rlabel metal2 s 52182 159200 52238 160800 6 reg_peri_rdata[14]
port 296 nsew signal input
rlabel metal2 s 51998 159200 52054 160800 6 reg_peri_rdata[15]
port 297 nsew signal input
rlabel metal2 s 51814 159200 51870 160800 6 reg_peri_rdata[16]
port 298 nsew signal input
rlabel metal2 s 51630 159200 51686 160800 6 reg_peri_rdata[17]
port 299 nsew signal input
rlabel metal2 s 51446 159200 51502 160800 6 reg_peri_rdata[18]
port 300 nsew signal input
rlabel metal2 s 51262 159200 51318 160800 6 reg_peri_rdata[19]
port 301 nsew signal input
rlabel metal2 s 54574 159200 54630 160800 6 reg_peri_rdata[1]
port 302 nsew signal input
rlabel metal2 s 51078 159200 51134 160800 6 reg_peri_rdata[20]
port 303 nsew signal input
rlabel metal2 s 50894 159200 50950 160800 6 reg_peri_rdata[21]
port 304 nsew signal input
rlabel metal2 s 50710 159200 50766 160800 6 reg_peri_rdata[22]
port 305 nsew signal input
rlabel metal2 s 50526 159200 50582 160800 6 reg_peri_rdata[23]
port 306 nsew signal input
rlabel metal2 s 50342 159200 50398 160800 6 reg_peri_rdata[24]
port 307 nsew signal input
rlabel metal2 s 50158 159200 50214 160800 6 reg_peri_rdata[25]
port 308 nsew signal input
rlabel metal2 s 49974 159200 50030 160800 6 reg_peri_rdata[26]
port 309 nsew signal input
rlabel metal2 s 49790 159200 49846 160800 6 reg_peri_rdata[27]
port 310 nsew signal input
rlabel metal2 s 49606 159200 49662 160800 6 reg_peri_rdata[28]
port 311 nsew signal input
rlabel metal2 s 49422 159200 49478 160800 6 reg_peri_rdata[29]
port 312 nsew signal input
rlabel metal2 s 54390 159200 54446 160800 6 reg_peri_rdata[2]
port 313 nsew signal input
rlabel metal2 s 49238 159200 49294 160800 6 reg_peri_rdata[30]
port 314 nsew signal input
rlabel metal2 s 49054 159200 49110 160800 6 reg_peri_rdata[31]
port 315 nsew signal input
rlabel metal2 s 54206 159200 54262 160800 6 reg_peri_rdata[3]
port 316 nsew signal input
rlabel metal2 s 54022 159200 54078 160800 6 reg_peri_rdata[4]
port 317 nsew signal input
rlabel metal2 s 53838 159200 53894 160800 6 reg_peri_rdata[5]
port 318 nsew signal input
rlabel metal2 s 53654 159200 53710 160800 6 reg_peri_rdata[6]
port 319 nsew signal input
rlabel metal2 s 53470 159200 53526 160800 6 reg_peri_rdata[7]
port 320 nsew signal input
rlabel metal2 s 53286 159200 53342 160800 6 reg_peri_rdata[8]
port 321 nsew signal input
rlabel metal2 s 53102 159200 53158 160800 6 reg_peri_rdata[9]
port 322 nsew signal input
rlabel metal2 s 48870 159200 48926 160800 6 reg_peri_wdata[0]
port 323 nsew signal output
rlabel metal2 s 47030 159200 47086 160800 6 reg_peri_wdata[10]
port 324 nsew signal output
rlabel metal2 s 46846 159200 46902 160800 6 reg_peri_wdata[11]
port 325 nsew signal output
rlabel metal2 s 46662 159200 46718 160800 6 reg_peri_wdata[12]
port 326 nsew signal output
rlabel metal2 s 46478 159200 46534 160800 6 reg_peri_wdata[13]
port 327 nsew signal output
rlabel metal2 s 46294 159200 46350 160800 6 reg_peri_wdata[14]
port 328 nsew signal output
rlabel metal2 s 46110 159200 46166 160800 6 reg_peri_wdata[15]
port 329 nsew signal output
rlabel metal2 s 45926 159200 45982 160800 6 reg_peri_wdata[16]
port 330 nsew signal output
rlabel metal2 s 45742 159200 45798 160800 6 reg_peri_wdata[17]
port 331 nsew signal output
rlabel metal2 s 45558 159200 45614 160800 6 reg_peri_wdata[18]
port 332 nsew signal output
rlabel metal2 s 45374 159200 45430 160800 6 reg_peri_wdata[19]
port 333 nsew signal output
rlabel metal2 s 48686 159200 48742 160800 6 reg_peri_wdata[1]
port 334 nsew signal output
rlabel metal2 s 45190 159200 45246 160800 6 reg_peri_wdata[20]
port 335 nsew signal output
rlabel metal2 s 45006 159200 45062 160800 6 reg_peri_wdata[21]
port 336 nsew signal output
rlabel metal2 s 44822 159200 44878 160800 6 reg_peri_wdata[22]
port 337 nsew signal output
rlabel metal2 s 44638 159200 44694 160800 6 reg_peri_wdata[23]
port 338 nsew signal output
rlabel metal2 s 44454 159200 44510 160800 6 reg_peri_wdata[24]
port 339 nsew signal output
rlabel metal2 s 44270 159200 44326 160800 6 reg_peri_wdata[25]
port 340 nsew signal output
rlabel metal2 s 44086 159200 44142 160800 6 reg_peri_wdata[26]
port 341 nsew signal output
rlabel metal2 s 43902 159200 43958 160800 6 reg_peri_wdata[27]
port 342 nsew signal output
rlabel metal2 s 43718 159200 43774 160800 6 reg_peri_wdata[28]
port 343 nsew signal output
rlabel metal2 s 43534 159200 43590 160800 6 reg_peri_wdata[29]
port 344 nsew signal output
rlabel metal2 s 48502 159200 48558 160800 6 reg_peri_wdata[2]
port 345 nsew signal output
rlabel metal2 s 43350 159200 43406 160800 6 reg_peri_wdata[30]
port 346 nsew signal output
rlabel metal2 s 43166 159200 43222 160800 6 reg_peri_wdata[31]
port 347 nsew signal output
rlabel metal2 s 48318 159200 48374 160800 6 reg_peri_wdata[3]
port 348 nsew signal output
rlabel metal2 s 48134 159200 48190 160800 6 reg_peri_wdata[4]
port 349 nsew signal output
rlabel metal2 s 47950 159200 48006 160800 6 reg_peri_wdata[5]
port 350 nsew signal output
rlabel metal2 s 47766 159200 47822 160800 6 reg_peri_wdata[6]
port 351 nsew signal output
rlabel metal2 s 47582 159200 47638 160800 6 reg_peri_wdata[7]
port 352 nsew signal output
rlabel metal2 s 47398 159200 47454 160800 6 reg_peri_wdata[8]
port 353 nsew signal output
rlabel metal2 s 47214 159200 47270 160800 6 reg_peri_wdata[9]
port 354 nsew signal output
rlabel metal2 s 40222 159200 40278 160800 6 reg_peri_wr
port 355 nsew signal output
rlabel metal3 s -800 73856 800 73976 4 reg_rdata[0]
port 356 nsew signal output
rlabel metal3 s -800 71136 800 71256 4 reg_rdata[10]
port 357 nsew signal output
rlabel metal3 s -800 70864 800 70984 4 reg_rdata[11]
port 358 nsew signal output
rlabel metal3 s -800 70592 800 70712 4 reg_rdata[12]
port 359 nsew signal output
rlabel metal3 s -800 70320 800 70440 4 reg_rdata[13]
port 360 nsew signal output
rlabel metal3 s -800 70048 800 70168 4 reg_rdata[14]
port 361 nsew signal output
rlabel metal3 s -800 69776 800 69896 4 reg_rdata[15]
port 362 nsew signal output
rlabel metal3 s -800 69504 800 69624 4 reg_rdata[16]
port 363 nsew signal output
rlabel metal3 s -800 69232 800 69352 4 reg_rdata[17]
port 364 nsew signal output
rlabel metal3 s -800 68960 800 69080 4 reg_rdata[18]
port 365 nsew signal output
rlabel metal3 s -800 68688 800 68808 4 reg_rdata[19]
port 366 nsew signal output
rlabel metal3 s -800 73584 800 73704 4 reg_rdata[1]
port 367 nsew signal output
rlabel metal3 s -800 68416 800 68536 4 reg_rdata[20]
port 368 nsew signal output
rlabel metal3 s -800 68144 800 68264 4 reg_rdata[21]
port 369 nsew signal output
rlabel metal3 s -800 67872 800 67992 4 reg_rdata[22]
port 370 nsew signal output
rlabel metal3 s -800 67600 800 67720 4 reg_rdata[23]
port 371 nsew signal output
rlabel metal3 s -800 67328 800 67448 4 reg_rdata[24]
port 372 nsew signal output
rlabel metal3 s -800 67056 800 67176 4 reg_rdata[25]
port 373 nsew signal output
rlabel metal3 s -800 66784 800 66904 4 reg_rdata[26]
port 374 nsew signal output
rlabel metal3 s -800 66512 800 66632 4 reg_rdata[27]
port 375 nsew signal output
rlabel metal3 s -800 66240 800 66360 4 reg_rdata[28]
port 376 nsew signal output
rlabel metal3 s -800 65968 800 66088 4 reg_rdata[29]
port 377 nsew signal output
rlabel metal3 s -800 73312 800 73432 4 reg_rdata[2]
port 378 nsew signal output
rlabel metal3 s -800 65696 800 65816 4 reg_rdata[30]
port 379 nsew signal output
rlabel metal3 s -800 65424 800 65544 4 reg_rdata[31]
port 380 nsew signal output
rlabel metal3 s -800 73040 800 73160 4 reg_rdata[3]
port 381 nsew signal output
rlabel metal3 s -800 72768 800 72888 4 reg_rdata[4]
port 382 nsew signal output
rlabel metal3 s -800 72496 800 72616 4 reg_rdata[5]
port 383 nsew signal output
rlabel metal3 s -800 72224 800 72344 4 reg_rdata[6]
port 384 nsew signal output
rlabel metal3 s -800 71952 800 72072 4 reg_rdata[7]
port 385 nsew signal output
rlabel metal3 s -800 71680 800 71800 4 reg_rdata[8]
port 386 nsew signal output
rlabel metal3 s -800 71408 800 71528 4 reg_rdata[9]
port 387 nsew signal output
rlabel metal3 s -800 65152 800 65272 4 reg_wdata[0]
port 388 nsew signal input
rlabel metal3 s -800 62432 800 62552 4 reg_wdata[10]
port 389 nsew signal input
rlabel metal3 s -800 62160 800 62280 4 reg_wdata[11]
port 390 nsew signal input
rlabel metal3 s -800 61888 800 62008 4 reg_wdata[12]
port 391 nsew signal input
rlabel metal3 s -800 61616 800 61736 4 reg_wdata[13]
port 392 nsew signal input
rlabel metal3 s -800 61344 800 61464 4 reg_wdata[14]
port 393 nsew signal input
rlabel metal3 s -800 61072 800 61192 4 reg_wdata[15]
port 394 nsew signal input
rlabel metal3 s -800 60800 800 60920 4 reg_wdata[16]
port 395 nsew signal input
rlabel metal3 s -800 60528 800 60648 4 reg_wdata[17]
port 396 nsew signal input
rlabel metal3 s -800 60256 800 60376 4 reg_wdata[18]
port 397 nsew signal input
rlabel metal3 s -800 59984 800 60104 4 reg_wdata[19]
port 398 nsew signal input
rlabel metal3 s -800 64880 800 65000 4 reg_wdata[1]
port 399 nsew signal input
rlabel metal3 s -800 59712 800 59832 4 reg_wdata[20]
port 400 nsew signal input
rlabel metal3 s -800 59440 800 59560 4 reg_wdata[21]
port 401 nsew signal input
rlabel metal3 s -800 59168 800 59288 4 reg_wdata[22]
port 402 nsew signal input
rlabel metal3 s -800 58896 800 59016 4 reg_wdata[23]
port 403 nsew signal input
rlabel metal3 s -800 58624 800 58744 4 reg_wdata[24]
port 404 nsew signal input
rlabel metal3 s -800 58352 800 58472 4 reg_wdata[25]
port 405 nsew signal input
rlabel metal3 s -800 58080 800 58200 4 reg_wdata[26]
port 406 nsew signal input
rlabel metal3 s -800 57808 800 57928 4 reg_wdata[27]
port 407 nsew signal input
rlabel metal3 s -800 57536 800 57656 4 reg_wdata[28]
port 408 nsew signal input
rlabel metal3 s -800 57264 800 57384 4 reg_wdata[29]
port 409 nsew signal input
rlabel metal3 s -800 64608 800 64728 4 reg_wdata[2]
port 410 nsew signal input
rlabel metal3 s -800 56992 800 57112 4 reg_wdata[30]
port 411 nsew signal input
rlabel metal3 s -800 56720 800 56840 4 reg_wdata[31]
port 412 nsew signal input
rlabel metal3 s -800 64336 800 64456 4 reg_wdata[3]
port 413 nsew signal input
rlabel metal3 s -800 64064 800 64184 4 reg_wdata[4]
port 414 nsew signal input
rlabel metal3 s -800 63792 800 63912 4 reg_wdata[5]
port 415 nsew signal input
rlabel metal3 s -800 63520 800 63640 4 reg_wdata[6]
port 416 nsew signal input
rlabel metal3 s -800 63248 800 63368 4 reg_wdata[7]
port 417 nsew signal input
rlabel metal3 s -800 62976 800 63096 4 reg_wdata[8]
port 418 nsew signal input
rlabel metal3 s -800 62704 800 62824 4 reg_wdata[9]
port 419 nsew signal input
rlabel metal3 s -800 52368 800 52488 4 reg_wr
port 420 nsew signal input
rlabel metal3 s -800 140360 800 140480 4 riscv_tck
port 421 nsew signal output
rlabel metal3 s -800 140904 800 141024 4 riscv_tdi
port 422 nsew signal output
rlabel metal3 s -800 141176 800 141296 4 riscv_tdo
port 423 nsew signal input
rlabel metal3 s -800 141448 800 141568 4 riscv_tdo_en
port 424 nsew signal input
rlabel metal3 s -800 140632 800 140752 4 riscv_tms
port 425 nsew signal output
rlabel metal3 s -800 140088 800 140208 4 riscv_trst_n
port 426 nsew signal output
rlabel metal2 s 30102 159200 30158 160800 6 rtc_clk
port 427 nsew signal output
rlabel metal2 s 30286 159200 30342 160800 6 rtc_intr
port 428 nsew signal input
rlabel metal2 s 21546 -800 21602 800 8 s_reset_n
port 429 nsew signal input
rlabel metal3 s 103200 3680 104800 3800 6 sflash_di[0]
port 430 nsew signal output
rlabel metal3 s 103200 3952 104800 4072 6 sflash_di[1]
port 431 nsew signal output
rlabel metal3 s 103200 4224 104800 4344 6 sflash_di[2]
port 432 nsew signal output
rlabel metal3 s 103200 4496 104800 4616 6 sflash_di[3]
port 433 nsew signal output
rlabel metal3 s 103200 2592 104800 2712 6 sflash_do[0]
port 434 nsew signal input
rlabel metal3 s 103200 2864 104800 2984 6 sflash_do[1]
port 435 nsew signal input
rlabel metal3 s 103200 3136 104800 3256 6 sflash_do[2]
port 436 nsew signal input
rlabel metal3 s 103200 3408 104800 3528 6 sflash_do[3]
port 437 nsew signal input
rlabel metal3 s 103200 144 104800 264 6 sflash_oen[0]
port 438 nsew signal input
rlabel metal3 s 103200 416 104800 536 6 sflash_oen[1]
port 439 nsew signal input
rlabel metal3 s 103200 688 104800 808 6 sflash_oen[2]
port 440 nsew signal input
rlabel metal3 s 103200 960 104800 1080 6 sflash_oen[3]
port 441 nsew signal input
rlabel metal3 s 103200 2320 104800 2440 6 sflash_sck
port 442 nsew signal input
rlabel metal3 s 103200 1232 104800 1352 6 sflash_ss[0]
port 443 nsew signal input
rlabel metal3 s 103200 1504 104800 1624 6 sflash_ss[1]
port 444 nsew signal input
rlabel metal3 s 103200 1776 104800 1896 6 sflash_ss[2]
port 445 nsew signal input
rlabel metal3 s 103200 2048 104800 2168 6 sflash_ss[3]
port 446 nsew signal input
rlabel metal2 s 31022 159200 31078 160800 6 sm_a1
port 447 nsew signal input
rlabel metal2 s 31206 159200 31262 160800 6 sm_a2
port 448 nsew signal input
rlabel metal2 s 31390 159200 31446 160800 6 sm_b1
port 449 nsew signal input
rlabel metal2 s 31574 159200 31630 160800 6 sm_b2
port 450 nsew signal input
rlabel metal3 s -800 40128 800 40248 4 soft_irq
port 451 nsew signal output
rlabel metal2 s 9310 -800 9366 800 8 spim_miso
port 452 nsew signal input
rlabel metal2 s 9494 -800 9550 800 8 spim_mosi
port 453 nsew signal output
rlabel metal2 s 8390 -800 8446 800 8 spim_sck
port 454 nsew signal input
rlabel metal2 s 9126 -800 9182 800 8 spim_ssn[0]
port 455 nsew signal input
rlabel metal2 s 8942 -800 8998 800 8 spim_ssn[1]
port 456 nsew signal input
rlabel metal2 s 8758 -800 8814 800 8 spim_ssn[2]
port 457 nsew signal input
rlabel metal2 s 8574 -800 8630 800 8 spim_ssn[3]
port 458 nsew signal input
rlabel metal2 s 10966 -800 11022 800 8 spis_miso
port 459 nsew signal input
rlabel metal2 s 11150 -800 11206 800 8 spis_mosi
port 460 nsew signal output
rlabel metal2 s 10598 -800 10654 800 8 spis_sck
port 461 nsew signal output
rlabel metal2 s 10782 -800 10838 800 8 spis_ssn
port 462 nsew signal output
rlabel metal2 s 1214 -800 1270 800 8 sspim_rst_n
port 463 nsew signal output
rlabel metal3 s -800 8576 800 8696 4 strap_sticky[0]
port 464 nsew signal output
rlabel metal3 s -800 5856 800 5976 4 strap_sticky[10]
port 465 nsew signal output
rlabel metal3 s -800 5584 800 5704 4 strap_sticky[11]
port 466 nsew signal output
rlabel metal3 s -800 5312 800 5432 4 strap_sticky[12]
port 467 nsew signal output
rlabel metal3 s -800 5040 800 5160 4 strap_sticky[13]
port 468 nsew signal output
rlabel metal3 s -800 4768 800 4888 4 strap_sticky[14]
port 469 nsew signal output
rlabel metal3 s -800 4496 800 4616 4 strap_sticky[15]
port 470 nsew signal output
rlabel metal3 s -800 4224 800 4344 4 strap_sticky[16]
port 471 nsew signal output
rlabel metal3 s -800 3952 800 4072 4 strap_sticky[17]
port 472 nsew signal output
rlabel metal3 s -800 3680 800 3800 4 strap_sticky[18]
port 473 nsew signal output
rlabel metal3 s -800 3408 800 3528 4 strap_sticky[19]
port 474 nsew signal output
rlabel metal3 s -800 8304 800 8424 4 strap_sticky[1]
port 475 nsew signal output
rlabel metal3 s -800 3136 800 3256 4 strap_sticky[20]
port 476 nsew signal output
rlabel metal3 s -800 2864 800 2984 4 strap_sticky[21]
port 477 nsew signal output
rlabel metal3 s -800 2592 800 2712 4 strap_sticky[22]
port 478 nsew signal output
rlabel metal3 s -800 2320 800 2440 4 strap_sticky[23]
port 479 nsew signal output
rlabel metal3 s -800 2048 800 2168 4 strap_sticky[24]
port 480 nsew signal output
rlabel metal3 s -800 1776 800 1896 4 strap_sticky[25]
port 481 nsew signal output
rlabel metal3 s -800 1504 800 1624 4 strap_sticky[26]
port 482 nsew signal output
rlabel metal3 s -800 1232 800 1352 4 strap_sticky[27]
port 483 nsew signal output
rlabel metal3 s -800 960 800 1080 4 strap_sticky[28]
port 484 nsew signal output
rlabel metal3 s -800 688 800 808 4 strap_sticky[29]
port 485 nsew signal output
rlabel metal3 s -800 8032 800 8152 4 strap_sticky[2]
port 486 nsew signal output
rlabel metal3 s -800 416 800 536 4 strap_sticky[30]
port 487 nsew signal output
rlabel metal3 s -800 144 800 264 4 strap_sticky[31]
port 488 nsew signal output
rlabel metal3 s -800 7760 800 7880 4 strap_sticky[3]
port 489 nsew signal output
rlabel metal3 s -800 7488 800 7608 4 strap_sticky[4]
port 490 nsew signal output
rlabel metal3 s -800 7216 800 7336 4 strap_sticky[5]
port 491 nsew signal output
rlabel metal3 s -800 6944 800 7064 4 strap_sticky[6]
port 492 nsew signal output
rlabel metal3 s -800 6672 800 6792 4 strap_sticky[7]
port 493 nsew signal output
rlabel metal3 s -800 6400 800 6520 4 strap_sticky[8]
port 494 nsew signal output
rlabel metal3 s -800 6128 800 6248 4 strap_sticky[9]
port 495 nsew signal output
rlabel metal3 s -800 9120 800 9240 4 strap_uartm[0]
port 496 nsew signal output
rlabel metal3 s -800 8848 800 8968 4 strap_uartm[1]
port 497 nsew signal output
rlabel metal3 s -800 17824 800 17944 4 system_strap[0]
port 498 nsew signal input
rlabel metal3 s -800 15104 800 15224 4 system_strap[10]
port 499 nsew signal input
rlabel metal3 s -800 14832 800 14952 4 system_strap[11]
port 500 nsew signal input
rlabel metal3 s -800 14560 800 14680 4 system_strap[12]
port 501 nsew signal input
rlabel metal3 s -800 14288 800 14408 4 system_strap[13]
port 502 nsew signal input
rlabel metal3 s -800 14016 800 14136 4 system_strap[14]
port 503 nsew signal input
rlabel metal3 s -800 13744 800 13864 4 system_strap[15]
port 504 nsew signal input
rlabel metal3 s -800 13472 800 13592 4 system_strap[16]
port 505 nsew signal input
rlabel metal3 s -800 13200 800 13320 4 system_strap[17]
port 506 nsew signal input
rlabel metal3 s -800 12928 800 13048 4 system_strap[18]
port 507 nsew signal input
rlabel metal3 s -800 12656 800 12776 4 system_strap[19]
port 508 nsew signal input
rlabel metal3 s -800 17552 800 17672 4 system_strap[1]
port 509 nsew signal input
rlabel metal3 s -800 12384 800 12504 4 system_strap[20]
port 510 nsew signal input
rlabel metal3 s -800 12112 800 12232 4 system_strap[21]
port 511 nsew signal input
rlabel metal3 s -800 11840 800 11960 4 system_strap[22]
port 512 nsew signal input
rlabel metal3 s -800 11568 800 11688 4 system_strap[23]
port 513 nsew signal input
rlabel metal3 s -800 11296 800 11416 4 system_strap[24]
port 514 nsew signal input
rlabel metal3 s -800 11024 800 11144 4 system_strap[25]
port 515 nsew signal input
rlabel metal3 s -800 10752 800 10872 4 system_strap[26]
port 516 nsew signal input
rlabel metal3 s -800 10480 800 10600 4 system_strap[27]
port 517 nsew signal input
rlabel metal3 s -800 10208 800 10328 4 system_strap[28]
port 518 nsew signal input
rlabel metal3 s -800 9936 800 10056 4 system_strap[29]
port 519 nsew signal input
rlabel metal3 s -800 17280 800 17400 4 system_strap[2]
port 520 nsew signal input
rlabel metal3 s -800 9664 800 9784 4 system_strap[30]
port 521 nsew signal input
rlabel metal3 s -800 9392 800 9512 4 system_strap[31]
port 522 nsew signal input
rlabel metal3 s -800 17008 800 17128 4 system_strap[3]
port 523 nsew signal input
rlabel metal3 s -800 16736 800 16856 4 system_strap[4]
port 524 nsew signal input
rlabel metal3 s -800 16464 800 16584 4 system_strap[5]
port 525 nsew signal input
rlabel metal3 s -800 16192 800 16312 4 system_strap[6]
port 526 nsew signal input
rlabel metal3 s -800 15920 800 16040 4 system_strap[7]
port 527 nsew signal input
rlabel metal3 s -800 15648 800 15768 4 system_strap[8]
port 528 nsew signal input
rlabel metal3 s -800 15376 800 15496 4 system_strap[9]
port 529 nsew signal input
rlabel metal2 s 1582 -800 1638 800 8 uart_rst_n[0]
port 530 nsew signal output
rlabel metal2 s 1398 -800 1454 800 8 uart_rst_n[1]
port 531 nsew signal output
rlabel metal2 s 7102 -800 7158 800 8 uart_rxd[0]
port 532 nsew signal output
rlabel metal2 s 6734 -800 6790 800 8 uart_rxd[1]
port 533 nsew signal output
rlabel metal2 s 6918 -800 6974 800 8 uart_txd[0]
port 534 nsew signal input
rlabel metal2 s 6550 -800 6606 800 8 uart_txd[1]
port 535 nsew signal input
rlabel metal2 s 10230 -800 10286 800 8 uartm_rxd
port 536 nsew signal output
rlabel metal2 s 10414 -800 10470 800 8 uartm_txd
port 537 nsew signal input
rlabel metal2 s 21914 -800 21970 800 8 usb_clk
port 538 nsew signal output
rlabel metal2 s 6366 -800 6422 800 8 usb_dn_i
port 539 nsew signal output
rlabel metal2 s 5814 -800 5870 800 8 usb_dn_o
port 540 nsew signal input
rlabel metal2 s 6182 -800 6238 800 8 usb_dp_i
port 541 nsew signal output
rlabel metal2 s 5630 -800 5686 800 8 usb_dp_o
port 542 nsew signal input
rlabel metal2 s 10046 -800 10102 800 8 usb_intr
port 543 nsew signal input
rlabel metal2 s 5998 -800 6054 800 8 usb_oen
port 544 nsew signal input
rlabel metal2 s 1950 -800 2006 800 8 usb_rst_n
port 545 nsew signal output
rlabel metal2 s 20074 -800 20130 800 8 user_clock1
port 546 nsew signal input
rlabel metal2 s 20442 -800 20498 800 8 user_clock2
port 547 nsew signal input
rlabel metal2 s 5078 -800 5134 800 8 user_irq[0]
port 548 nsew signal output
rlabel metal2 s 5262 -800 5318 800 8 user_irq[1]
port 549 nsew signal output
rlabel metal2 s 5446 -800 5502 800 8 user_irq[2]
port 550 nsew signal output
rlabel metal4 s 3748 2128 4988 157808 6 vccd1
port 551 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 157808 6 vccd1
port 551 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 157808 6 vccd1
port 551 nsew power bidirectional
rlabel metal4 s 63748 2128 64988 157808 6 vccd1
port 551 nsew power bidirectional
rlabel metal4 s 83748 2128 84988 157808 6 vccd1
port 551 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 157808 6 vssd1
port 552 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 157808 6 vssd1
port 552 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 157808 6 vssd1
port 552 nsew ground bidirectional
rlabel metal4 s 73748 2128 74988 157808 6 vssd1
port 552 nsew ground bidirectional
rlabel metal4 s 93748 2128 94988 157808 6 vssd1
port 552 nsew ground bidirectional
rlabel metal3 s -800 50192 800 50312 4 wbd_clk_int
port 553 nsew signal input
rlabel metal3 s -800 50464 800 50584 4 wbd_clk_pinmux
port 554 nsew signal output
rlabel metal2 s 21178 -800 21234 800 8 xtal_clk
port 555 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 104000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 49588312
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/pinmux_top/runs/pinmux_top/results/signoff/pinmux_top.magic.gds
string GDS_START 1336244
<< end >>

