magic
tech sky130A
magscale 1 2
timestamp 1698814312
<< obsli1 >>
rect 1104 2159 58880 357425
<< obsm1 >>
rect 14 348 59970 357456
<< metal2 >>
rect 110 0 166 800
rect 294 0 350 800
rect 478 0 534 800
rect 4066 0 4122 800
rect 4250 0 4306 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5170 0 5226 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 6090 0 6146 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 7010 0 7066 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7930 0 7986 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8850 0 8906 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9770 0 9826 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10690 0 10746 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11610 0 11666 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12530 0 12586 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 13082 0 13138 800
rect 13266 0 13322 800
rect 13450 0 13506 800
rect 13634 0 13690 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20442 0 20498 800
rect 20626 0 20682 800
rect 20810 0 20866 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21362 0 21418 800
rect 21546 0 21602 800
rect 21730 0 21786 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22282 0 22338 800
rect 22466 0 22522 800
rect 22650 0 22706 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23202 0 23258 800
rect 23386 0 23442 800
rect 23570 0 23626 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24122 0 24178 800
rect 24306 0 24362 800
rect 24490 0 24546 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 25042 0 25098 800
rect 25226 0 25282 800
rect 25410 0 25466 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25962 0 26018 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26882 0 26938 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27802 0 27858 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28722 0 28778 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29642 0 29698 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30562 0 30618 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31482 0 31538 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32402 0 32458 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33322 0 33378 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34242 0 34298 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35162 0 35218 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 36082 0 36138 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 37002 0 37058 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37922 0 37978 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38842 0 38898 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39394 0 39450 800
rect 45098 0 45154 800
rect 45282 0 45338 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45834 0 45890 800
rect 46018 0 46074 800
rect 46202 0 46258 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46754 0 46810 800
rect 46938 0 46994 800
rect 47122 0 47178 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47674 0 47730 800
rect 47858 0 47914 800
rect 48042 0 48098 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48594 0 48650 800
rect 48778 0 48834 800
rect 48962 0 49018 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49514 0 49570 800
rect 49698 0 49754 800
rect 49882 0 49938 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50434 0 50490 800
rect 50618 0 50674 800
rect 50802 0 50858 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51354 0 51410 800
rect 51538 0 51594 800
rect 51722 0 51778 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52274 0 52330 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53194 0 53250 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54114 0 54170 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 55034 0 55090 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55954 0 56010 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56874 0 56930 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57794 0 57850 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58714 0 58770 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59634 0 59690 800
rect 59818 0 59874 800
<< obsm2 >>
rect 20 856 59964 357445
rect 20 167 54 856
rect 222 167 238 856
rect 406 167 422 856
rect 590 167 4010 856
rect 4178 167 4194 856
rect 4362 167 4378 856
rect 4546 167 4562 856
rect 4730 167 4746 856
rect 4914 167 4930 856
rect 5098 167 5114 856
rect 5282 167 5298 856
rect 5466 167 5482 856
rect 5650 167 5666 856
rect 5834 167 5850 856
rect 6018 167 6034 856
rect 6202 167 6218 856
rect 6386 167 6402 856
rect 6570 167 6586 856
rect 6754 167 6770 856
rect 6938 167 6954 856
rect 7122 167 7138 856
rect 7306 167 7322 856
rect 7490 167 7506 856
rect 7674 167 7690 856
rect 7858 167 7874 856
rect 8042 167 8058 856
rect 8226 167 8242 856
rect 8410 167 8426 856
rect 8594 167 8610 856
rect 8778 167 8794 856
rect 8962 167 8978 856
rect 9146 167 9162 856
rect 9330 167 9346 856
rect 9514 167 9530 856
rect 9698 167 9714 856
rect 9882 167 9898 856
rect 10066 167 10082 856
rect 10250 167 10266 856
rect 10434 167 10450 856
rect 10618 167 10634 856
rect 10802 167 10818 856
rect 10986 167 11002 856
rect 11170 167 11186 856
rect 11354 167 11370 856
rect 11538 167 11554 856
rect 11722 167 11738 856
rect 11906 167 11922 856
rect 12090 167 12106 856
rect 12274 167 12290 856
rect 12458 167 12474 856
rect 12642 167 12658 856
rect 12826 167 12842 856
rect 13010 167 13026 856
rect 13194 167 13210 856
rect 13378 167 13394 856
rect 13562 167 13578 856
rect 13746 167 20018 856
rect 20186 167 20202 856
rect 20370 167 20386 856
rect 20554 167 20570 856
rect 20738 167 20754 856
rect 20922 167 20938 856
rect 21106 167 21122 856
rect 21290 167 21306 856
rect 21474 167 21490 856
rect 21658 167 21674 856
rect 21842 167 21858 856
rect 22026 167 22042 856
rect 22210 167 22226 856
rect 22394 167 22410 856
rect 22578 167 22594 856
rect 22762 167 22778 856
rect 22946 167 22962 856
rect 23130 167 23146 856
rect 23314 167 23330 856
rect 23498 167 23514 856
rect 23682 167 23698 856
rect 23866 167 23882 856
rect 24050 167 24066 856
rect 24234 167 24250 856
rect 24418 167 24434 856
rect 24602 167 24618 856
rect 24786 167 24802 856
rect 24970 167 24986 856
rect 25154 167 25170 856
rect 25338 167 25354 856
rect 25522 167 25538 856
rect 25706 167 25722 856
rect 25890 167 25906 856
rect 26074 167 26090 856
rect 26258 167 26274 856
rect 26442 167 26458 856
rect 26626 167 26642 856
rect 26810 167 26826 856
rect 26994 167 27010 856
rect 27178 167 27194 856
rect 27362 167 27378 856
rect 27546 167 27562 856
rect 27730 167 27746 856
rect 27914 167 27930 856
rect 28098 167 28114 856
rect 28282 167 28298 856
rect 28466 167 28482 856
rect 28650 167 28666 856
rect 28834 167 28850 856
rect 29018 167 29034 856
rect 29202 167 29218 856
rect 29386 167 29402 856
rect 29570 167 29586 856
rect 29754 167 29770 856
rect 29938 167 29954 856
rect 30122 167 30138 856
rect 30306 167 30322 856
rect 30490 167 30506 856
rect 30674 167 30690 856
rect 30858 167 30874 856
rect 31042 167 31058 856
rect 31226 167 31242 856
rect 31410 167 31426 856
rect 31594 167 31610 856
rect 31778 167 31794 856
rect 31962 167 31978 856
rect 32146 167 32162 856
rect 32330 167 32346 856
rect 32514 167 32530 856
rect 32698 167 32714 856
rect 32882 167 32898 856
rect 33066 167 33082 856
rect 33250 167 33266 856
rect 33434 167 33450 856
rect 33618 167 33634 856
rect 33802 167 33818 856
rect 33986 167 34002 856
rect 34170 167 34186 856
rect 34354 167 34370 856
rect 34538 167 34554 856
rect 34722 167 34738 856
rect 34906 167 34922 856
rect 35090 167 35106 856
rect 35274 167 35290 856
rect 35458 167 35474 856
rect 35642 167 35658 856
rect 35826 167 35842 856
rect 36010 167 36026 856
rect 36194 167 36210 856
rect 36378 167 36394 856
rect 36562 167 36578 856
rect 36746 167 36762 856
rect 36930 167 36946 856
rect 37114 167 37130 856
rect 37298 167 37314 856
rect 37482 167 37498 856
rect 37666 167 37682 856
rect 37850 167 37866 856
rect 38034 167 38050 856
rect 38218 167 38234 856
rect 38402 167 38418 856
rect 38586 167 38602 856
rect 38770 167 38786 856
rect 38954 167 38970 856
rect 39138 167 39154 856
rect 39322 167 39338 856
rect 39506 167 45042 856
rect 45210 167 45226 856
rect 45394 167 45410 856
rect 45578 167 45594 856
rect 45762 167 45778 856
rect 45946 167 45962 856
rect 46130 167 46146 856
rect 46314 167 46330 856
rect 46498 167 46514 856
rect 46682 167 46698 856
rect 46866 167 46882 856
rect 47050 167 47066 856
rect 47234 167 47250 856
rect 47418 167 47434 856
rect 47602 167 47618 856
rect 47786 167 47802 856
rect 47970 167 47986 856
rect 48154 167 48170 856
rect 48338 167 48354 856
rect 48522 167 48538 856
rect 48706 167 48722 856
rect 48890 167 48906 856
rect 49074 167 49090 856
rect 49258 167 49274 856
rect 49442 167 49458 856
rect 49626 167 49642 856
rect 49810 167 49826 856
rect 49994 167 50010 856
rect 50178 167 50194 856
rect 50362 167 50378 856
rect 50546 167 50562 856
rect 50730 167 50746 856
rect 50914 167 50930 856
rect 51098 167 51114 856
rect 51282 167 51298 856
rect 51466 167 51482 856
rect 51650 167 51666 856
rect 51834 167 51850 856
rect 52018 167 52034 856
rect 52202 167 52218 856
rect 52386 167 52402 856
rect 52570 167 52586 856
rect 52754 167 52770 856
rect 52938 167 52954 856
rect 53122 167 53138 856
rect 53306 167 53322 856
rect 53490 167 53506 856
rect 53674 167 53690 856
rect 53858 167 53874 856
rect 54042 167 54058 856
rect 54226 167 54242 856
rect 54410 167 54426 856
rect 54594 167 54610 856
rect 54778 167 54794 856
rect 54962 167 54978 856
rect 55146 167 55162 856
rect 55330 167 55346 856
rect 55514 167 55530 856
rect 55698 167 55714 856
rect 55882 167 55898 856
rect 56066 167 56082 856
rect 56250 167 56266 856
rect 56434 167 56450 856
rect 56618 167 56634 856
rect 56802 167 56818 856
rect 56986 167 57002 856
rect 57170 167 57186 856
rect 57354 167 57370 856
rect 57538 167 57554 856
rect 57722 167 57738 856
rect 57906 167 57922 856
rect 58090 167 58106 856
rect 58274 167 58290 856
rect 58458 167 58474 856
rect 58642 167 58658 856
rect 58826 167 58842 856
rect 59010 167 59026 856
rect 59194 167 59210 856
rect 59378 167 59394 856
rect 59562 167 59578 856
rect 59746 167 59762 856
rect 59930 167 59964 856
<< metal3 >>
rect 59200 351160 60000 351280
rect 0 350888 800 351008
rect 0 350616 800 350736
rect 0 350344 800 350464
rect 0 350072 800 350192
rect 59200 350888 60000 351008
rect 59200 350616 60000 350736
rect 59200 350344 60000 350464
rect 59200 350072 60000 350192
rect 0 340960 800 341080
rect 0 340688 800 340808
rect 0 340416 800 340536
rect 0 340144 800 340264
rect 0 328720 800 328840
rect 0 328448 800 328568
rect 0 328176 800 328296
rect 0 327904 800 328024
rect 0 327632 800 327752
rect 0 327360 800 327480
rect 0 327088 800 327208
rect 0 326816 800 326936
rect 0 326544 800 326664
rect 0 326272 800 326392
rect 0 326000 800 326120
rect 0 325728 800 325848
rect 0 325456 800 325576
rect 0 325184 800 325304
rect 0 324912 800 325032
rect 0 324640 800 324760
rect 0 324368 800 324488
rect 0 324096 800 324216
rect 0 323824 800 323944
rect 0 323552 800 323672
rect 0 323280 800 323400
rect 0 323008 800 323128
rect 0 322736 800 322856
rect 0 322464 800 322584
rect 0 322192 800 322312
rect 0 321920 800 322040
rect 0 321648 800 321768
rect 0 321376 800 321496
rect 0 321104 800 321224
rect 0 320832 800 320952
rect 0 320560 800 320680
rect 0 320288 800 320408
rect 0 320016 800 320136
rect 59200 304648 60000 304768
rect 59200 304376 60000 304496
rect 59200 304104 60000 304224
rect 59200 303832 60000 303952
rect 59200 303560 60000 303680
rect 59200 303288 60000 303408
rect 59200 303016 60000 303136
rect 59200 302744 60000 302864
rect 59200 302472 60000 302592
rect 59200 302200 60000 302320
rect 59200 301928 60000 302048
rect 59200 301656 60000 301776
rect 59200 301384 60000 301504
rect 59200 301112 60000 301232
rect 59200 300840 60000 300960
rect 59200 300568 60000 300688
rect 59200 300296 60000 300416
rect 59200 300024 60000 300144
rect 59200 299752 60000 299872
rect 59200 299480 60000 299600
rect 59200 299208 60000 299328
rect 59200 298936 60000 299056
rect 59200 298664 60000 298784
rect 59200 298392 60000 298512
rect 59200 298120 60000 298240
rect 59200 297848 60000 297968
rect 59200 297576 60000 297696
rect 59200 297304 60000 297424
rect 59200 297032 60000 297152
rect 59200 296760 60000 296880
rect 59200 296488 60000 296608
rect 59200 296216 60000 296336
rect 59200 295944 60000 296064
rect 59200 295672 60000 295792
rect 59200 295400 60000 295520
rect 59200 295128 60000 295248
rect 59200 294856 60000 294976
rect 59200 294584 60000 294704
rect 59200 294312 60000 294432
rect 59200 294040 60000 294160
rect 59200 293768 60000 293888
rect 59200 293496 60000 293616
rect 59200 293224 60000 293344
rect 59200 292952 60000 293072
rect 59200 292680 60000 292800
rect 59200 292408 60000 292528
rect 59200 292136 60000 292256
rect 59200 291864 60000 291984
rect 59200 291592 60000 291712
rect 59200 291320 60000 291440
rect 59200 291048 60000 291168
rect 59200 290776 60000 290896
rect 59200 290504 60000 290624
rect 59200 290232 60000 290352
rect 59200 289960 60000 290080
rect 59200 289688 60000 289808
rect 59200 289416 60000 289536
rect 59200 289144 60000 289264
rect 59200 288872 60000 288992
rect 59200 288600 60000 288720
rect 59200 288328 60000 288448
rect 59200 288056 60000 288176
rect 59200 287784 60000 287904
rect 59200 287512 60000 287632
rect 59200 287240 60000 287360
rect 59200 286968 60000 287088
rect 59200 286696 60000 286816
rect 59200 286424 60000 286544
rect 59200 286152 60000 286272
rect 59200 285880 60000 286000
rect 59200 285608 60000 285728
rect 59200 285336 60000 285456
rect 59200 285064 60000 285184
rect 59200 284792 60000 284912
rect 59200 284520 60000 284640
rect 59200 284248 60000 284368
rect 59200 283976 60000 284096
rect 59200 283704 60000 283824
rect 59200 283432 60000 283552
rect 59200 283160 60000 283280
rect 59200 282888 60000 283008
rect 59200 282616 60000 282736
rect 59200 282344 60000 282464
rect 59200 282072 60000 282192
rect 59200 279896 60000 280016
rect 59200 279624 60000 279744
rect 59200 279352 60000 279472
rect 59200 279080 60000 279200
rect 59200 278808 60000 278928
rect 59200 278536 60000 278656
rect 59200 278264 60000 278384
rect 59200 277992 60000 278112
rect 59200 277720 60000 277840
rect 59200 277448 60000 277568
rect 59200 277176 60000 277296
rect 59200 276904 60000 277024
rect 59200 276632 60000 276752
rect 59200 276360 60000 276480
rect 59200 276088 60000 276208
rect 59200 275816 60000 275936
rect 59200 275544 60000 275664
rect 59200 275272 60000 275392
rect 59200 275000 60000 275120
rect 59200 274728 60000 274848
rect 59200 274456 60000 274576
rect 59200 274184 60000 274304
rect 59200 273912 60000 274032
rect 59200 273640 60000 273760
rect 59200 273368 60000 273488
rect 59200 273096 60000 273216
rect 59200 272824 60000 272944
rect 59200 272552 60000 272672
rect 59200 272280 60000 272400
rect 59200 272008 60000 272128
rect 59200 271736 60000 271856
rect 59200 271464 60000 271584
rect 59200 271192 60000 271312
rect 59200 270920 60000 271040
rect 59200 270648 60000 270768
rect 59200 270376 60000 270496
rect 59200 270104 60000 270224
rect 59200 248616 60000 248736
rect 59200 248344 60000 248464
rect 59200 248072 60000 248192
rect 59200 247800 60000 247920
rect 59200 247528 60000 247648
rect 59200 247256 60000 247376
rect 59200 246984 60000 247104
rect 59200 246712 60000 246832
rect 59200 246440 60000 246560
rect 59200 246168 60000 246288
rect 59200 245896 60000 246016
rect 59200 245624 60000 245744
rect 59200 245352 60000 245472
rect 59200 245080 60000 245200
rect 59200 244808 60000 244928
rect 59200 244536 60000 244656
rect 59200 244264 60000 244384
rect 59200 243992 60000 244112
rect 59200 243720 60000 243840
rect 59200 243448 60000 243568
rect 59200 243176 60000 243296
rect 59200 242904 60000 243024
rect 59200 242632 60000 242752
rect 59200 242360 60000 242480
rect 59200 242088 60000 242208
rect 59200 241816 60000 241936
rect 59200 241544 60000 241664
rect 59200 241272 60000 241392
rect 59200 241000 60000 241120
rect 59200 240728 60000 240848
rect 59200 240456 60000 240576
rect 59200 240184 60000 240304
rect 59200 239912 60000 240032
rect 59200 239640 60000 239760
rect 59200 239368 60000 239488
rect 59200 239096 60000 239216
rect 59200 238824 60000 238944
rect 59200 238552 60000 238672
rect 59200 238280 60000 238400
rect 59200 238008 60000 238128
rect 59200 237736 60000 237856
rect 59200 237464 60000 237584
rect 59200 237192 60000 237312
rect 59200 236920 60000 237040
rect 59200 236648 60000 236768
rect 59200 236376 60000 236496
rect 59200 236104 60000 236224
rect 59200 235832 60000 235952
rect 59200 235560 60000 235680
rect 59200 235288 60000 235408
rect 59200 235016 60000 235136
rect 59200 234744 60000 234864
rect 59200 234472 60000 234592
rect 59200 234200 60000 234320
rect 59200 233928 60000 234048
rect 59200 233656 60000 233776
rect 59200 233384 60000 233504
rect 59200 233112 60000 233232
rect 59200 232840 60000 232960
rect 59200 232568 60000 232688
rect 59200 232296 60000 232416
rect 59200 232024 60000 232144
rect 59200 231752 60000 231872
rect 59200 231480 60000 231600
rect 59200 231208 60000 231328
rect 59200 230936 60000 231056
rect 59200 230664 60000 230784
rect 59200 230392 60000 230512
rect 59200 230120 60000 230240
rect 59200 172048 60000 172168
rect 59200 171776 60000 171896
rect 59200 171504 60000 171624
rect 59200 171232 60000 171352
rect 59200 170960 60000 171080
rect 59200 170688 60000 170808
rect 59200 170416 60000 170536
rect 59200 170144 60000 170264
rect 59200 169872 60000 169992
rect 59200 169600 60000 169720
rect 59200 169328 60000 169448
rect 59200 169056 60000 169176
rect 59200 168784 60000 168904
rect 59200 168512 60000 168632
rect 59200 168240 60000 168360
rect 59200 167968 60000 168088
rect 59200 167696 60000 167816
rect 59200 167424 60000 167544
rect 59200 167152 60000 167272
rect 59200 166880 60000 167000
rect 59200 166608 60000 166728
rect 59200 166336 60000 166456
rect 59200 166064 60000 166184
rect 59200 165792 60000 165912
rect 59200 165520 60000 165640
rect 59200 165248 60000 165368
rect 59200 164976 60000 165096
rect 59200 164704 60000 164824
rect 59200 164432 60000 164552
rect 59200 164160 60000 164280
rect 59200 163888 60000 164008
rect 59200 163616 60000 163736
rect 59200 163344 60000 163464
rect 59200 163072 60000 163192
rect 59200 162800 60000 162920
rect 59200 162528 60000 162648
rect 59200 162256 60000 162376
rect 59200 161984 60000 162104
rect 59200 161712 60000 161832
rect 59200 161440 60000 161560
rect 59200 161168 60000 161288
rect 59200 160896 60000 161016
rect 59200 160624 60000 160744
rect 59200 160352 60000 160472
rect 59200 160080 60000 160200
rect 59200 159808 60000 159928
rect 59200 159536 60000 159656
rect 59200 159264 60000 159384
rect 59200 158992 60000 159112
rect 59200 158720 60000 158840
rect 59200 158448 60000 158568
rect 59200 158176 60000 158296
rect 59200 157904 60000 158024
rect 59200 157632 60000 157752
rect 59200 157360 60000 157480
rect 59200 157088 60000 157208
rect 59200 156816 60000 156936
rect 59200 156544 60000 156664
rect 59200 156272 60000 156392
rect 59200 156000 60000 156120
rect 59200 155728 60000 155848
rect 59200 155456 60000 155576
rect 59200 155184 60000 155304
rect 59200 154912 60000 155032
rect 59200 154640 60000 154760
rect 59200 154368 60000 154488
rect 59200 154096 60000 154216
rect 59200 153824 60000 153944
rect 59200 153552 60000 153672
rect 59200 153280 60000 153400
rect 59200 153008 60000 153128
rect 59200 152736 60000 152856
rect 59200 152464 60000 152584
rect 59200 152192 60000 152312
rect 59200 151920 60000 152040
rect 59200 151648 60000 151768
rect 59200 151376 60000 151496
rect 0 151104 800 151224
rect 0 150832 800 150952
rect 0 150560 800 150680
rect 0 150288 800 150408
rect 0 150016 800 150136
rect 59200 151104 60000 151224
rect 59200 150832 60000 150952
rect 59200 150560 60000 150680
rect 59200 150288 60000 150408
rect 59200 150016 60000 150136
rect 0 134376 800 134496
rect 0 134104 800 134224
rect 0 133832 800 133952
rect 0 133560 800 133680
rect 0 133288 800 133408
rect 0 133016 800 133136
rect 0 132744 800 132864
rect 0 132472 800 132592
rect 0 132200 800 132320
rect 0 131928 800 132048
rect 0 131656 800 131776
rect 0 131384 800 131504
rect 0 131112 800 131232
rect 0 130840 800 130960
rect 0 130568 800 130688
rect 0 130296 800 130416
rect 0 130024 800 130144
rect 59200 130840 60000 130960
rect 59200 130568 60000 130688
rect 59200 130296 60000 130416
rect 59200 130024 60000 130144
rect 0 122952 800 123072
rect 0 122680 800 122800
rect 0 122408 800 122528
rect 0 122136 800 122256
rect 0 121864 800 121984
rect 0 121592 800 121712
rect 0 121320 800 121440
rect 0 121048 800 121168
rect 0 120776 800 120896
rect 0 120504 800 120624
rect 0 120232 800 120352
rect 0 119960 800 120080
rect 0 119688 800 119808
rect 0 119416 800 119536
rect 0 119144 800 119264
rect 0 118872 800 118992
rect 0 118600 800 118720
rect 0 118328 800 118448
rect 0 118056 800 118176
rect 0 117784 800 117904
rect 0 117512 800 117632
rect 0 117240 800 117360
rect 0 116968 800 117088
rect 0 116696 800 116816
rect 0 116424 800 116544
rect 0 116152 800 116272
rect 0 115880 800 116000
rect 0 115608 800 115728
rect 0 115336 800 115456
rect 0 115064 800 115184
rect 0 114792 800 114912
rect 0 114520 800 114640
rect 0 114248 800 114368
rect 0 113976 800 114096
rect 0 113704 800 113824
rect 0 113432 800 113552
rect 0 113160 800 113280
rect 0 112888 800 113008
rect 0 112616 800 112736
rect 0 112344 800 112464
rect 0 112072 800 112192
rect 0 111800 800 111920
rect 0 111528 800 111648
rect 0 111256 800 111376
rect 0 110984 800 111104
rect 0 110712 800 110832
rect 0 110440 800 110560
rect 0 110168 800 110288
rect 0 109896 800 110016
rect 0 109624 800 109744
rect 0 109352 800 109472
rect 0 109080 800 109200
rect 0 108808 800 108928
rect 0 108536 800 108656
rect 0 108264 800 108384
rect 0 107992 800 108112
rect 0 107720 800 107840
rect 0 107448 800 107568
rect 0 107176 800 107296
rect 0 106904 800 107024
rect 0 106632 800 106752
rect 0 106360 800 106480
rect 0 106088 800 106208
rect 0 105816 800 105936
rect 0 105544 800 105664
rect 0 105272 800 105392
rect 0 105000 800 105120
rect 0 104728 800 104848
rect 0 104456 800 104576
rect 0 104184 800 104304
rect 0 103912 800 104032
rect 0 103640 800 103760
rect 0 103368 800 103488
rect 0 103096 800 103216
rect 0 102824 800 102944
rect 0 102552 800 102672
rect 0 102280 800 102400
rect 0 102008 800 102128
rect 0 101736 800 101856
rect 0 101464 800 101584
rect 0 101192 800 101312
rect 0 100920 800 101040
rect 0 100648 800 100768
rect 0 100376 800 100496
rect 0 100104 800 100224
rect 0 91672 800 91792
rect 0 91400 800 91520
rect 0 91128 800 91248
rect 0 90856 800 90976
rect 0 90584 800 90704
rect 0 90312 800 90432
rect 0 90040 800 90160
rect 0 89768 800 89888
rect 0 89496 800 89616
rect 0 89224 800 89344
rect 0 88952 800 89072
rect 0 88680 800 88800
rect 0 88408 800 88528
rect 0 88136 800 88256
rect 0 87864 800 87984
rect 0 87592 800 87712
rect 0 87320 800 87440
rect 0 87048 800 87168
rect 0 86776 800 86896
rect 0 86504 800 86624
rect 0 86232 800 86352
rect 0 85960 800 86080
rect 0 85688 800 85808
rect 0 85416 800 85536
rect 0 85144 800 85264
rect 0 84872 800 84992
rect 0 84600 800 84720
rect 0 84328 800 84448
rect 0 84056 800 84176
rect 0 83784 800 83904
rect 0 83512 800 83632
rect 0 83240 800 83360
rect 0 82968 800 83088
rect 0 82696 800 82816
rect 0 82424 800 82544
rect 0 82152 800 82272
rect 0 81880 800 82000
rect 0 81608 800 81728
rect 0 81336 800 81456
rect 0 81064 800 81184
rect 0 80792 800 80912
rect 0 80520 800 80640
rect 0 80248 800 80368
rect 0 79976 800 80096
rect 0 79704 800 79824
rect 0 79432 800 79552
rect 0 79160 800 79280
rect 0 78888 800 79008
rect 0 78616 800 78736
rect 0 78344 800 78464
rect 0 78072 800 78192
rect 0 77800 800 77920
rect 0 77528 800 77648
rect 0 77256 800 77376
rect 0 76984 800 77104
rect 0 76712 800 76832
rect 0 76440 800 76560
rect 0 76168 800 76288
rect 0 75896 800 76016
rect 0 75624 800 75744
rect 0 75352 800 75472
rect 0 75080 800 75200
rect 0 74808 800 74928
rect 0 74536 800 74656
rect 0 74264 800 74384
rect 0 73992 800 74112
rect 0 73720 800 73840
rect 0 73448 800 73568
rect 0 73176 800 73296
rect 0 72904 800 73024
rect 0 72632 800 72752
rect 0 72360 800 72480
rect 0 72088 800 72208
rect 0 71816 800 71936
rect 0 71544 800 71664
rect 0 71272 800 71392
rect 0 71000 800 71120
rect 0 70728 800 70848
rect 0 70456 800 70576
rect 0 70184 800 70304
rect 0 69912 800 70032
rect 0 69640 800 69760
rect 0 69368 800 69488
rect 0 69096 800 69216
rect 0 68824 800 68944
rect 0 68552 800 68672
rect 0 68280 800 68400
rect 0 68008 800 68128
rect 0 67736 800 67856
rect 0 67464 800 67584
rect 0 67192 800 67312
rect 0 66920 800 67040
rect 0 66648 800 66768
rect 0 66376 800 66496
rect 0 66104 800 66224
rect 0 65832 800 65952
rect 0 65560 800 65680
rect 0 65288 800 65408
rect 0 65016 800 65136
rect 0 64744 800 64864
rect 0 64472 800 64592
rect 0 64200 800 64320
rect 0 63928 800 64048
rect 0 63656 800 63776
rect 0 63384 800 63504
rect 0 63112 800 63232
rect 0 62840 800 62960
rect 0 62568 800 62688
rect 0 62296 800 62416
rect 0 62024 800 62144
rect 0 61752 800 61872
rect 0 61480 800 61600
rect 0 61208 800 61328
rect 0 60936 800 61056
rect 0 60664 800 60784
rect 0 60392 800 60512
rect 0 60120 800 60240
rect 0 49784 800 49904
rect 0 49512 800 49632
rect 0 49240 800 49360
rect 0 48968 800 49088
rect 0 48696 800 48816
rect 0 48424 800 48544
rect 0 48152 800 48272
rect 0 47880 800 48000
rect 0 47608 800 47728
rect 0 47336 800 47456
rect 0 47064 800 47184
rect 0 46792 800 46912
rect 0 46520 800 46640
rect 0 46248 800 46368
rect 0 45976 800 46096
rect 0 45704 800 45824
rect 0 45432 800 45552
rect 0 45160 800 45280
rect 0 44888 800 45008
rect 0 44616 800 44736
rect 0 44344 800 44464
rect 0 44072 800 44192
rect 0 43800 800 43920
rect 0 43528 800 43648
rect 0 43256 800 43376
rect 0 42984 800 43104
rect 0 42712 800 42832
rect 0 42440 800 42560
rect 0 42168 800 42288
rect 0 41896 800 42016
rect 0 41624 800 41744
rect 0 41352 800 41472
rect 0 41080 800 41200
rect 0 40808 800 40928
rect 0 40536 800 40656
rect 0 40264 800 40384
rect 0 39992 800 40112
rect 0 39720 800 39840
rect 0 39448 800 39568
rect 0 39176 800 39296
rect 0 38904 800 39024
rect 0 38632 800 38752
rect 0 38360 800 38480
rect 0 38088 800 38208
rect 0 37816 800 37936
rect 0 37544 800 37664
rect 0 37272 800 37392
rect 0 37000 800 37120
rect 0 36728 800 36848
rect 0 36456 800 36576
rect 0 36184 800 36304
rect 0 35912 800 36032
rect 0 35640 800 35760
rect 0 35368 800 35488
rect 0 35096 800 35216
rect 0 34824 800 34944
rect 0 34552 800 34672
rect 0 34280 800 34400
rect 0 34008 800 34128
rect 0 33736 800 33856
rect 0 33464 800 33584
rect 0 33192 800 33312
rect 0 32920 800 33040
rect 0 32648 800 32768
rect 0 32376 800 32496
rect 0 32104 800 32224
rect 0 31832 800 31952
rect 0 31560 800 31680
rect 0 31288 800 31408
rect 0 31016 800 31136
rect 0 30744 800 30864
rect 0 30472 800 30592
rect 0 30200 800 30320
rect 0 29928 800 30048
rect 0 29656 800 29776
rect 0 29384 800 29504
rect 0 29112 800 29232
rect 0 28840 800 28960
rect 0 28568 800 28688
rect 0 28296 800 28416
rect 0 28024 800 28144
rect 0 27752 800 27872
rect 0 27480 800 27600
rect 0 27208 800 27328
rect 0 26936 800 27056
rect 0 26664 800 26784
rect 0 26392 800 26512
rect 0 26120 800 26240
rect 0 25848 800 25968
rect 0 25576 800 25696
rect 0 25304 800 25424
rect 0 25032 800 25152
rect 0 24760 800 24880
rect 0 24488 800 24608
rect 0 24216 800 24336
rect 0 23944 800 24064
rect 0 23672 800 23792
rect 0 23400 800 23520
rect 0 23128 800 23248
rect 0 22856 800 22976
rect 0 22584 800 22704
rect 0 22312 800 22432
rect 0 22040 800 22160
rect 0 21768 800 21888
rect 0 21496 800 21616
rect 0 21224 800 21344
rect 0 20952 800 21072
rect 0 20680 800 20800
rect 0 20408 800 20528
rect 0 20136 800 20256
rect 59200 41896 60000 42016
rect 59200 41624 60000 41744
rect 59200 41352 60000 41472
rect 59200 41080 60000 41200
rect 59200 40808 60000 40928
rect 59200 40536 60000 40656
rect 59200 40264 60000 40384
rect 59200 39992 60000 40112
rect 59200 39720 60000 39840
rect 59200 39448 60000 39568
rect 59200 39176 60000 39296
rect 59200 38904 60000 39024
rect 59200 38632 60000 38752
rect 59200 38360 60000 38480
rect 59200 38088 60000 38208
rect 59200 37816 60000 37936
rect 59200 37544 60000 37664
rect 59200 37272 60000 37392
rect 59200 37000 60000 37120
rect 59200 36728 60000 36848
rect 59200 36456 60000 36576
rect 59200 36184 60000 36304
rect 59200 35912 60000 36032
rect 59200 35640 60000 35760
rect 59200 35368 60000 35488
rect 59200 35096 60000 35216
rect 59200 34824 60000 34944
rect 59200 34552 60000 34672
rect 59200 34280 60000 34400
rect 59200 34008 60000 34128
rect 59200 33736 60000 33856
rect 59200 33464 60000 33584
rect 59200 33192 60000 33312
rect 59200 32920 60000 33040
rect 59200 32648 60000 32768
rect 59200 32376 60000 32496
rect 59200 32104 60000 32224
rect 59200 31832 60000 31952
rect 59200 31560 60000 31680
rect 59200 31288 60000 31408
rect 59200 31016 60000 31136
rect 59200 30744 60000 30864
rect 59200 30472 60000 30592
rect 59200 30200 60000 30320
rect 59200 29928 60000 30048
rect 59200 29656 60000 29776
rect 59200 29384 60000 29504
rect 59200 29112 60000 29232
rect 59200 28840 60000 28960
rect 59200 28568 60000 28688
rect 59200 28296 60000 28416
rect 59200 28024 60000 28144
rect 59200 27752 60000 27872
rect 59200 27480 60000 27600
rect 59200 27208 60000 27328
rect 59200 26936 60000 27056
rect 59200 26664 60000 26784
rect 59200 26392 60000 26512
rect 59200 26120 60000 26240
rect 59200 25848 60000 25968
rect 59200 25576 60000 25696
rect 59200 25304 60000 25424
rect 59200 25032 60000 25152
rect 59200 24760 60000 24880
rect 59200 24488 60000 24608
rect 59200 24216 60000 24336
rect 59200 23944 60000 24064
rect 59200 23672 60000 23792
rect 59200 23400 60000 23520
rect 59200 23128 60000 23248
rect 59200 22856 60000 22976
rect 59200 22584 60000 22704
rect 59200 22312 60000 22432
rect 59200 22040 60000 22160
rect 59200 21768 60000 21888
rect 59200 21496 60000 21616
rect 59200 21224 60000 21344
rect 59200 20952 60000 21072
rect 59200 20680 60000 20800
rect 59200 20408 60000 20528
rect 59200 20136 60000 20256
rect 59200 19864 60000 19984
rect 59200 19592 60000 19712
rect 59200 19320 60000 19440
rect 59200 19048 60000 19168
rect 59200 18776 60000 18896
rect 59200 18504 60000 18624
rect 59200 18232 60000 18352
rect 59200 17960 60000 18080
rect 59200 17688 60000 17808
rect 59200 17416 60000 17536
rect 59200 17144 60000 17264
rect 59200 16872 60000 16992
rect 59200 16600 60000 16720
rect 59200 16328 60000 16448
rect 59200 16056 60000 16176
rect 59200 15784 60000 15904
rect 59200 15512 60000 15632
rect 59200 15240 60000 15360
rect 59200 14968 60000 15088
rect 59200 14696 60000 14816
rect 59200 14424 60000 14544
rect 59200 14152 60000 14272
rect 59200 13880 60000 14000
rect 59200 13608 60000 13728
rect 59200 13336 60000 13456
rect 59200 13064 60000 13184
rect 59200 12792 60000 12912
rect 59200 12520 60000 12640
rect 59200 12248 60000 12368
rect 59200 11976 60000 12096
rect 59200 11704 60000 11824
rect 59200 11432 60000 11552
rect 0 11160 800 11280
rect 0 10888 800 11008
rect 0 10616 800 10736
rect 0 10344 800 10464
rect 0 10072 800 10192
rect 59200 11160 60000 11280
rect 59200 10888 60000 11008
rect 59200 10616 60000 10736
rect 59200 10344 60000 10464
rect 59200 10072 60000 10192
rect 59200 2048 60000 2168
rect 59200 1776 60000 1896
rect 59200 1504 60000 1624
rect 0 1232 800 1352
rect 0 960 800 1080
rect 0 688 800 808
rect 0 416 800 536
rect 0 144 800 264
rect 59200 1232 60000 1352
rect 59200 960 60000 1080
rect 59200 688 60000 808
rect 59200 416 60000 536
rect 59200 144 60000 264
<< obsm3 >>
rect 54 351360 59235 357441
rect 54 351088 59120 351360
rect 880 349992 59120 351088
rect 54 341160 59235 349992
rect 880 340064 59235 341160
rect 54 328920 59235 340064
rect 880 319936 59235 328920
rect 54 304848 59235 319936
rect 54 281992 59120 304848
rect 54 280096 59235 281992
rect 54 270024 59120 280096
rect 54 248816 59235 270024
rect 54 230040 59120 248816
rect 54 172248 59235 230040
rect 54 151304 59120 172248
rect 880 149936 59120 151304
rect 54 134576 59235 149936
rect 880 131040 59235 134576
rect 880 129944 59120 131040
rect 54 123152 59235 129944
rect 880 100024 59235 123152
rect 54 91872 59235 100024
rect 880 60040 59235 91872
rect 54 49984 59235 60040
rect 880 42096 59235 49984
rect 880 20056 59120 42096
rect 54 11360 59120 20056
rect 880 9992 59120 11360
rect 54 2248 59235 9992
rect 54 1432 59120 2248
rect 880 171 59120 1432
<< metal4 >>
rect 3748 2128 4988 357456
rect 13748 2128 14988 357456
rect 23748 2128 24988 357456
rect 33748 2128 34988 357456
rect 43748 2128 44988 357456
rect 53748 2128 54988 357456
<< obsm4 >>
rect 59 2483 3668 350709
rect 5068 2483 13668 350709
rect 15068 2483 23668 350709
rect 25068 2483 33668 350709
rect 35068 2483 43668 350709
rect 45068 2483 53668 350709
rect 55068 2483 59005 350709
<< labels >>
rlabel metal2 s 12898 0 12954 800 6 cfg_cska_wi[0]
port 1 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 cfg_cska_wi[1]
port 2 nsew signal input
rlabel metal2 s 12530 0 12586 800 6 cfg_cska_wi[2]
port 3 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 cfg_cska_wi[3]
port 4 nsew signal input
rlabel metal2 s 478 0 534 800 6 ch_clk_in[0]
port 5 nsew signal input
rlabel metal2 s 294 0 350 800 6 ch_clk_in[1]
port 6 nsew signal input
rlabel metal2 s 110 0 166 800 6 ch_clk_in[2]
port 7 nsew signal input
rlabel metal3 s 0 1232 800 1352 6 ch_clk_out[0]
port 8 nsew signal output
rlabel metal3 s 0 134376 800 134496 6 ch_clk_out[1]
port 9 nsew signal output
rlabel metal3 s 0 151104 800 151224 6 ch_clk_out[2]
port 10 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 ch_data_in[0]
port 11 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 ch_data_in[100]
port 12 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 ch_data_in[101]
port 13 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 ch_data_in[102]
port 14 nsew signal input
rlabel metal2 s 55034 0 55090 800 6 ch_data_in[103]
port 15 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 ch_data_in[104]
port 16 nsew signal input
rlabel metal2 s 54666 0 54722 800 6 ch_data_in[105]
port 17 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 ch_data_in[106]
port 18 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 ch_data_in[107]
port 19 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 ch_data_in[108]
port 20 nsew signal input
rlabel metal2 s 53930 0 53986 800 6 ch_data_in[109]
port 21 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 ch_data_in[10]
port 22 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 ch_data_in[110]
port 23 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 ch_data_in[111]
port 24 nsew signal input
rlabel metal3 s 59200 239096 60000 239216 6 ch_data_in[112]
port 25 nsew signal input
rlabel metal3 s 59200 238824 60000 238944 6 ch_data_in[113]
port 26 nsew signal input
rlabel metal3 s 59200 238552 60000 238672 6 ch_data_in[114]
port 27 nsew signal input
rlabel metal3 s 59200 238280 60000 238400 6 ch_data_in[115]
port 28 nsew signal input
rlabel metal3 s 59200 238008 60000 238128 6 ch_data_in[116]
port 29 nsew signal input
rlabel metal3 s 59200 237736 60000 237856 6 ch_data_in[117]
port 30 nsew signal input
rlabel metal3 s 59200 237464 60000 237584 6 ch_data_in[118]
port 31 nsew signal input
rlabel metal3 s 59200 237192 60000 237312 6 ch_data_in[119]
port 32 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 ch_data_in[11]
port 33 nsew signal input
rlabel metal3 s 59200 236920 60000 237040 6 ch_data_in[120]
port 34 nsew signal input
rlabel metal3 s 59200 236648 60000 236768 6 ch_data_in[121]
port 35 nsew signal input
rlabel metal3 s 59200 236376 60000 236496 6 ch_data_in[122]
port 36 nsew signal input
rlabel metal3 s 59200 236104 60000 236224 6 ch_data_in[123]
port 37 nsew signal input
rlabel metal3 s 59200 235832 60000 235952 6 ch_data_in[124]
port 38 nsew signal input
rlabel metal3 s 59200 235560 60000 235680 6 ch_data_in[125]
port 39 nsew signal input
rlabel metal3 s 59200 235288 60000 235408 6 ch_data_in[126]
port 40 nsew signal input
rlabel metal3 s 59200 235016 60000 235136 6 ch_data_in[127]
port 41 nsew signal input
rlabel metal3 s 59200 234744 60000 234864 6 ch_data_in[128]
port 42 nsew signal input
rlabel metal3 s 59200 234472 60000 234592 6 ch_data_in[129]
port 43 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 ch_data_in[12]
port 44 nsew signal input
rlabel metal3 s 59200 234200 60000 234320 6 ch_data_in[130]
port 45 nsew signal input
rlabel metal3 s 59200 233928 60000 234048 6 ch_data_in[131]
port 46 nsew signal input
rlabel metal3 s 59200 233656 60000 233776 6 ch_data_in[132]
port 47 nsew signal input
rlabel metal3 s 59200 233384 60000 233504 6 ch_data_in[133]
port 48 nsew signal input
rlabel metal3 s 59200 233112 60000 233232 6 ch_data_in[134]
port 49 nsew signal input
rlabel metal3 s 59200 232840 60000 232960 6 ch_data_in[135]
port 50 nsew signal input
rlabel metal3 s 59200 232568 60000 232688 6 ch_data_in[136]
port 51 nsew signal input
rlabel metal3 s 59200 232296 60000 232416 6 ch_data_in[137]
port 52 nsew signal input
rlabel metal3 s 59200 232024 60000 232144 6 ch_data_in[138]
port 53 nsew signal input
rlabel metal3 s 59200 231752 60000 231872 6 ch_data_in[139]
port 54 nsew signal input
rlabel metal2 s 9770 0 9826 800 6 ch_data_in[13]
port 55 nsew signal input
rlabel metal3 s 59200 231480 60000 231600 6 ch_data_in[140]
port 56 nsew signal input
rlabel metal3 s 59200 231208 60000 231328 6 ch_data_in[141]
port 57 nsew signal input
rlabel metal3 s 59200 230936 60000 231056 6 ch_data_in[142]
port 58 nsew signal input
rlabel metal3 s 59200 230664 60000 230784 6 ch_data_in[143]
port 59 nsew signal input
rlabel metal3 s 59200 230392 60000 230512 6 ch_data_in[144]
port 60 nsew signal input
rlabel metal3 s 59200 230120 60000 230240 6 ch_data_in[145]
port 61 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 ch_data_in[146]
port 62 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 ch_data_in[147]
port 63 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 ch_data_in[148]
port 64 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 ch_data_in[149]
port 65 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 ch_data_in[14]
port 66 nsew signal input
rlabel metal2 s 46386 0 46442 800 6 ch_data_in[150]
port 67 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 ch_data_in[151]
port 68 nsew signal input
rlabel metal2 s 46018 0 46074 800 6 ch_data_in[152]
port 69 nsew signal input
rlabel metal2 s 45834 0 45890 800 6 ch_data_in[153]
port 70 nsew signal input
rlabel metal2 s 45650 0 45706 800 6 ch_data_in[154]
port 71 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 ch_data_in[155]
port 72 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 ch_data_in[156]
port 73 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 ch_data_in[157]
port 74 nsew signal input
rlabel metal2 s 9402 0 9458 800 6 ch_data_in[15]
port 75 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 ch_data_in[16]
port 76 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 ch_data_in[17]
port 77 nsew signal input
rlabel metal2 s 8850 0 8906 800 6 ch_data_in[18]
port 78 nsew signal input
rlabel metal2 s 8666 0 8722 800 6 ch_data_in[19]
port 79 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 ch_data_in[1]
port 80 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 ch_data_in[20]
port 81 nsew signal input
rlabel metal2 s 8298 0 8354 800 6 ch_data_in[21]
port 82 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 ch_data_in[22]
port 83 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 ch_data_in[23]
port 84 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 ch_data_in[24]
port 85 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 ch_data_in[25]
port 86 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 ch_data_in[26]
port 87 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 ch_data_in[27]
port 88 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 ch_data_in[28]
port 89 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 ch_data_in[29]
port 90 nsew signal input
rlabel metal2 s 11794 0 11850 800 6 ch_data_in[2]
port 91 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 ch_data_in[30]
port 92 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 ch_data_in[31]
port 93 nsew signal input
rlabel metal2 s 6274 0 6330 800 6 ch_data_in[32]
port 94 nsew signal input
rlabel metal2 s 6090 0 6146 800 6 ch_data_in[33]
port 95 nsew signal input
rlabel metal2 s 5906 0 5962 800 6 ch_data_in[34]
port 96 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 ch_data_in[35]
port 97 nsew signal input
rlabel metal2 s 5538 0 5594 800 6 ch_data_in[36]
port 98 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 ch_data_in[37]
port 99 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 ch_data_in[38]
port 100 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 ch_data_in[39]
port 101 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 ch_data_in[3]
port 102 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 ch_data_in[40]
port 103 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 ch_data_in[41]
port 104 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 ch_data_in[42]
port 105 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 ch_data_in[43]
port 106 nsew signal input
rlabel metal3 s 59200 278808 60000 278928 6 ch_data_in[44]
port 107 nsew signal input
rlabel metal3 s 59200 278536 60000 278656 6 ch_data_in[45]
port 108 nsew signal input
rlabel metal3 s 59200 278264 60000 278384 6 ch_data_in[46]
port 109 nsew signal input
rlabel metal3 s 59200 277992 60000 278112 6 ch_data_in[47]
port 110 nsew signal input
rlabel metal3 s 59200 277720 60000 277840 6 ch_data_in[48]
port 111 nsew signal input
rlabel metal3 s 59200 277448 60000 277568 6 ch_data_in[49]
port 112 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 ch_data_in[4]
port 113 nsew signal input
rlabel metal3 s 59200 277176 60000 277296 6 ch_data_in[50]
port 114 nsew signal input
rlabel metal3 s 59200 276904 60000 277024 6 ch_data_in[51]
port 115 nsew signal input
rlabel metal3 s 59200 276632 60000 276752 6 ch_data_in[52]
port 116 nsew signal input
rlabel metal3 s 59200 276360 60000 276480 6 ch_data_in[53]
port 117 nsew signal input
rlabel metal3 s 59200 276088 60000 276208 6 ch_data_in[54]
port 118 nsew signal input
rlabel metal3 s 59200 275816 60000 275936 6 ch_data_in[55]
port 119 nsew signal input
rlabel metal3 s 59200 275544 60000 275664 6 ch_data_in[56]
port 120 nsew signal input
rlabel metal3 s 59200 275272 60000 275392 6 ch_data_in[57]
port 121 nsew signal input
rlabel metal3 s 59200 275000 60000 275120 6 ch_data_in[58]
port 122 nsew signal input
rlabel metal3 s 59200 274728 60000 274848 6 ch_data_in[59]
port 123 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 ch_data_in[5]
port 124 nsew signal input
rlabel metal3 s 59200 274456 60000 274576 6 ch_data_in[60]
port 125 nsew signal input
rlabel metal3 s 59200 274184 60000 274304 6 ch_data_in[61]
port 126 nsew signal input
rlabel metal3 s 59200 273912 60000 274032 6 ch_data_in[62]
port 127 nsew signal input
rlabel metal3 s 59200 273640 60000 273760 6 ch_data_in[63]
port 128 nsew signal input
rlabel metal3 s 59200 273368 60000 273488 6 ch_data_in[64]
port 129 nsew signal input
rlabel metal3 s 59200 273096 60000 273216 6 ch_data_in[65]
port 130 nsew signal input
rlabel metal3 s 59200 272824 60000 272944 6 ch_data_in[66]
port 131 nsew signal input
rlabel metal3 s 59200 272552 60000 272672 6 ch_data_in[67]
port 132 nsew signal input
rlabel metal3 s 59200 272280 60000 272400 6 ch_data_in[68]
port 133 nsew signal input
rlabel metal3 s 59200 272008 60000 272128 6 ch_data_in[69]
port 134 nsew signal input
rlabel metal2 s 11058 0 11114 800 6 ch_data_in[6]
port 135 nsew signal input
rlabel metal3 s 59200 271736 60000 271856 6 ch_data_in[70]
port 136 nsew signal input
rlabel metal3 s 59200 271464 60000 271584 6 ch_data_in[71]
port 137 nsew signal input
rlabel metal3 s 59200 271192 60000 271312 6 ch_data_in[72]
port 138 nsew signal input
rlabel metal3 s 59200 270920 60000 271040 6 ch_data_in[73]
port 139 nsew signal input
rlabel metal3 s 59200 270648 60000 270768 6 ch_data_in[74]
port 140 nsew signal input
rlabel metal3 s 59200 270376 60000 270496 6 ch_data_in[75]
port 141 nsew signal input
rlabel metal3 s 59200 270104 60000 270224 6 ch_data_in[76]
port 142 nsew signal input
rlabel metal2 s 59818 0 59874 800 6 ch_data_in[77]
port 143 nsew signal input
rlabel metal2 s 59634 0 59690 800 6 ch_data_in[78]
port 144 nsew signal input
rlabel metal2 s 59450 0 59506 800 6 ch_data_in[79]
port 145 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 ch_data_in[7]
port 146 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 ch_data_in[80]
port 147 nsew signal input
rlabel metal2 s 59082 0 59138 800 6 ch_data_in[81]
port 148 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 ch_data_in[82]
port 149 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 ch_data_in[83]
port 150 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 ch_data_in[84]
port 151 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 ch_data_in[85]
port 152 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 ch_data_in[86]
port 153 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 ch_data_in[87]
port 154 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 ch_data_in[88]
port 155 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 ch_data_in[89]
port 156 nsew signal input
rlabel metal2 s 10690 0 10746 800 6 ch_data_in[8]
port 157 nsew signal input
rlabel metal2 s 57426 0 57482 800 6 ch_data_in[90]
port 158 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 ch_data_in[91]
port 159 nsew signal input
rlabel metal2 s 57058 0 57114 800 6 ch_data_in[92]
port 160 nsew signal input
rlabel metal2 s 56874 0 56930 800 6 ch_data_in[93]
port 161 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 ch_data_in[94]
port 162 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 ch_data_in[95]
port 163 nsew signal input
rlabel metal2 s 56322 0 56378 800 6 ch_data_in[96]
port 164 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 ch_data_in[97]
port 165 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 ch_data_in[98]
port 166 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 ch_data_in[99]
port 167 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 ch_data_in[9]
port 168 nsew signal input
rlabel metal3 s 0 10888 800 11008 6 ch_data_out[0]
port 169 nsew signal output
rlabel metal3 s 59200 242360 60000 242480 6 ch_data_out[100]
port 170 nsew signal output
rlabel metal3 s 59200 242088 60000 242208 6 ch_data_out[101]
port 171 nsew signal output
rlabel metal3 s 59200 241816 60000 241936 6 ch_data_out[102]
port 172 nsew signal output
rlabel metal3 s 59200 241544 60000 241664 6 ch_data_out[103]
port 173 nsew signal output
rlabel metal3 s 59200 241272 60000 241392 6 ch_data_out[104]
port 174 nsew signal output
rlabel metal3 s 59200 241000 60000 241120 6 ch_data_out[105]
port 175 nsew signal output
rlabel metal3 s 59200 240728 60000 240848 6 ch_data_out[106]
port 176 nsew signal output
rlabel metal3 s 59200 240456 60000 240576 6 ch_data_out[107]
port 177 nsew signal output
rlabel metal3 s 59200 240184 60000 240304 6 ch_data_out[108]
port 178 nsew signal output
rlabel metal3 s 59200 239912 60000 240032 6 ch_data_out[109]
port 179 nsew signal output
rlabel metal3 s 59200 130296 60000 130416 6 ch_data_out[10]
port 180 nsew signal output
rlabel metal3 s 59200 239640 60000 239760 6 ch_data_out[110]
port 181 nsew signal output
rlabel metal3 s 59200 239368 60000 239488 6 ch_data_out[111]
port 182 nsew signal output
rlabel metal2 s 53378 0 53434 800 6 ch_data_out[112]
port 183 nsew signal output
rlabel metal2 s 53194 0 53250 800 6 ch_data_out[113]
port 184 nsew signal output
rlabel metal2 s 53010 0 53066 800 6 ch_data_out[114]
port 185 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 ch_data_out[115]
port 186 nsew signal output
rlabel metal2 s 52642 0 52698 800 6 ch_data_out[116]
port 187 nsew signal output
rlabel metal2 s 52458 0 52514 800 6 ch_data_out[117]
port 188 nsew signal output
rlabel metal2 s 52274 0 52330 800 6 ch_data_out[118]
port 189 nsew signal output
rlabel metal2 s 52090 0 52146 800 6 ch_data_out[119]
port 190 nsew signal output
rlabel metal3 s 59200 130024 60000 130144 6 ch_data_out[11]
port 191 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 ch_data_out[120]
port 192 nsew signal output
rlabel metal2 s 51722 0 51778 800 6 ch_data_out[121]
port 193 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 ch_data_out[122]
port 194 nsew signal output
rlabel metal2 s 51354 0 51410 800 6 ch_data_out[123]
port 195 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 ch_data_out[124]
port 196 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 ch_data_out[125]
port 197 nsew signal output
rlabel metal2 s 50802 0 50858 800 6 ch_data_out[126]
port 198 nsew signal output
rlabel metal2 s 50618 0 50674 800 6 ch_data_out[127]
port 199 nsew signal output
rlabel metal2 s 50434 0 50490 800 6 ch_data_out[128]
port 200 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 ch_data_out[129]
port 201 nsew signal output
rlabel metal3 s 59200 279896 60000 280016 6 ch_data_out[12]
port 202 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 ch_data_out[130]
port 203 nsew signal output
rlabel metal2 s 49882 0 49938 800 6 ch_data_out[131]
port 204 nsew signal output
rlabel metal2 s 49698 0 49754 800 6 ch_data_out[132]
port 205 nsew signal output
rlabel metal2 s 49514 0 49570 800 6 ch_data_out[133]
port 206 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 ch_data_out[134]
port 207 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 ch_data_out[135]
port 208 nsew signal output
rlabel metal2 s 48962 0 49018 800 6 ch_data_out[136]
port 209 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 ch_data_out[137]
port 210 nsew signal output
rlabel metal2 s 48594 0 48650 800 6 ch_data_out[138]
port 211 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 ch_data_out[139]
port 212 nsew signal output
rlabel metal3 s 59200 279624 60000 279744 6 ch_data_out[13]
port 213 nsew signal output
rlabel metal2 s 48226 0 48282 800 6 ch_data_out[140]
port 214 nsew signal output
rlabel metal2 s 48042 0 48098 800 6 ch_data_out[141]
port 215 nsew signal output
rlabel metal2 s 47858 0 47914 800 6 ch_data_out[142]
port 216 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 ch_data_out[143]
port 217 nsew signal output
rlabel metal2 s 47490 0 47546 800 6 ch_data_out[144]
port 218 nsew signal output
rlabel metal2 s 47306 0 47362 800 6 ch_data_out[145]
port 219 nsew signal output
rlabel metal3 s 0 340960 800 341080 6 ch_data_out[146]
port 220 nsew signal output
rlabel metal3 s 0 340688 800 340808 6 ch_data_out[147]
port 221 nsew signal output
rlabel metal3 s 0 340416 800 340536 6 ch_data_out[148]
port 222 nsew signal output
rlabel metal3 s 0 340144 800 340264 6 ch_data_out[149]
port 223 nsew signal output
rlabel metal3 s 59200 279352 60000 279472 6 ch_data_out[14]
port 224 nsew signal output
rlabel metal3 s 0 350888 800 351008 6 ch_data_out[150]
port 225 nsew signal output
rlabel metal3 s 0 350616 800 350736 6 ch_data_out[151]
port 226 nsew signal output
rlabel metal3 s 0 350344 800 350464 6 ch_data_out[152]
port 227 nsew signal output
rlabel metal3 s 0 350072 800 350192 6 ch_data_out[153]
port 228 nsew signal output
rlabel metal3 s 59200 350344 60000 350464 6 ch_data_out[154]
port 229 nsew signal output
rlabel metal3 s 59200 350616 60000 350736 6 ch_data_out[155]
port 230 nsew signal output
rlabel metal3 s 59200 350888 60000 351008 6 ch_data_out[156]
port 231 nsew signal output
rlabel metal3 s 59200 351160 60000 351280 6 ch_data_out[157]
port 232 nsew signal output
rlabel metal3 s 59200 279080 60000 279200 6 ch_data_out[15]
port 233 nsew signal output
rlabel metal3 s 59200 960 60000 1080 6 ch_data_out[16]
port 234 nsew signal output
rlabel metal3 s 59200 688 60000 808 6 ch_data_out[17]
port 235 nsew signal output
rlabel metal3 s 59200 416 60000 536 6 ch_data_out[18]
port 236 nsew signal output
rlabel metal3 s 59200 144 60000 264 6 ch_data_out[19]
port 237 nsew signal output
rlabel metal3 s 0 10616 800 10736 6 ch_data_out[1]
port 238 nsew signal output
rlabel metal3 s 0 960 800 1080 6 ch_data_out[20]
port 239 nsew signal output
rlabel metal3 s 0 688 800 808 6 ch_data_out[21]
port 240 nsew signal output
rlabel metal3 s 0 416 800 536 6 ch_data_out[22]
port 241 nsew signal output
rlabel metal3 s 0 144 800 264 6 ch_data_out[23]
port 242 nsew signal output
rlabel metal3 s 0 150832 800 150952 6 ch_data_out[24]
port 243 nsew signal output
rlabel metal3 s 0 150560 800 150680 6 ch_data_out[25]
port 244 nsew signal output
rlabel metal3 s 0 150288 800 150408 6 ch_data_out[26]
port 245 nsew signal output
rlabel metal3 s 0 150016 800 150136 6 ch_data_out[27]
port 246 nsew signal output
rlabel metal3 s 0 134104 800 134224 6 ch_data_out[28]
port 247 nsew signal output
rlabel metal3 s 0 133832 800 133952 6 ch_data_out[29]
port 248 nsew signal output
rlabel metal3 s 0 10344 800 10464 6 ch_data_out[2]
port 249 nsew signal output
rlabel metal3 s 0 133560 800 133680 6 ch_data_out[30]
port 250 nsew signal output
rlabel metal3 s 0 133288 800 133408 6 ch_data_out[31]
port 251 nsew signal output
rlabel metal3 s 0 133016 800 133136 6 ch_data_out[32]
port 252 nsew signal output
rlabel metal3 s 0 132744 800 132864 6 ch_data_out[33]
port 253 nsew signal output
rlabel metal3 s 0 132472 800 132592 6 ch_data_out[34]
port 254 nsew signal output
rlabel metal3 s 0 132200 800 132320 6 ch_data_out[35]
port 255 nsew signal output
rlabel metal3 s 0 131928 800 132048 6 ch_data_out[36]
port 256 nsew signal output
rlabel metal3 s 0 131656 800 131776 6 ch_data_out[37]
port 257 nsew signal output
rlabel metal3 s 0 131384 800 131504 6 ch_data_out[38]
port 258 nsew signal output
rlabel metal3 s 0 131112 800 131232 6 ch_data_out[39]
port 259 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 ch_data_out[3]
port 260 nsew signal output
rlabel metal3 s 0 130840 800 130960 6 ch_data_out[40]
port 261 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 ch_data_out[41]
port 262 nsew signal output
rlabel metal3 s 0 130296 800 130416 6 ch_data_out[42]
port 263 nsew signal output
rlabel metal3 s 0 130024 800 130144 6 ch_data_out[43]
port 264 nsew signal output
rlabel metal3 s 0 328720 800 328840 6 ch_data_out[44]
port 265 nsew signal output
rlabel metal3 s 0 328448 800 328568 6 ch_data_out[45]
port 266 nsew signal output
rlabel metal3 s 0 328176 800 328296 6 ch_data_out[46]
port 267 nsew signal output
rlabel metal3 s 0 327904 800 328024 6 ch_data_out[47]
port 268 nsew signal output
rlabel metal3 s 0 327632 800 327752 6 ch_data_out[48]
port 269 nsew signal output
rlabel metal3 s 0 327360 800 327480 6 ch_data_out[49]
port 270 nsew signal output
rlabel metal3 s 59200 2048 60000 2168 6 ch_data_out[4]
port 271 nsew signal output
rlabel metal3 s 0 327088 800 327208 6 ch_data_out[50]
port 272 nsew signal output
rlabel metal3 s 0 326816 800 326936 6 ch_data_out[51]
port 273 nsew signal output
rlabel metal3 s 0 326544 800 326664 6 ch_data_out[52]
port 274 nsew signal output
rlabel metal3 s 0 326272 800 326392 6 ch_data_out[53]
port 275 nsew signal output
rlabel metal3 s 0 326000 800 326120 6 ch_data_out[54]
port 276 nsew signal output
rlabel metal3 s 0 325728 800 325848 6 ch_data_out[55]
port 277 nsew signal output
rlabel metal3 s 0 325456 800 325576 6 ch_data_out[56]
port 278 nsew signal output
rlabel metal3 s 0 325184 800 325304 6 ch_data_out[57]
port 279 nsew signal output
rlabel metal3 s 0 324912 800 325032 6 ch_data_out[58]
port 280 nsew signal output
rlabel metal3 s 0 324640 800 324760 6 ch_data_out[59]
port 281 nsew signal output
rlabel metal3 s 59200 1776 60000 1896 6 ch_data_out[5]
port 282 nsew signal output
rlabel metal3 s 0 324368 800 324488 6 ch_data_out[60]
port 283 nsew signal output
rlabel metal3 s 0 324096 800 324216 6 ch_data_out[61]
port 284 nsew signal output
rlabel metal3 s 0 323824 800 323944 6 ch_data_out[62]
port 285 nsew signal output
rlabel metal3 s 0 323552 800 323672 6 ch_data_out[63]
port 286 nsew signal output
rlabel metal3 s 0 323280 800 323400 6 ch_data_out[64]
port 287 nsew signal output
rlabel metal3 s 0 323008 800 323128 6 ch_data_out[65]
port 288 nsew signal output
rlabel metal3 s 0 322736 800 322856 6 ch_data_out[66]
port 289 nsew signal output
rlabel metal3 s 0 322464 800 322584 6 ch_data_out[67]
port 290 nsew signal output
rlabel metal3 s 0 322192 800 322312 6 ch_data_out[68]
port 291 nsew signal output
rlabel metal3 s 0 321920 800 322040 6 ch_data_out[69]
port 292 nsew signal output
rlabel metal3 s 59200 1504 60000 1624 6 ch_data_out[6]
port 293 nsew signal output
rlabel metal3 s 0 321648 800 321768 6 ch_data_out[70]
port 294 nsew signal output
rlabel metal3 s 0 321376 800 321496 6 ch_data_out[71]
port 295 nsew signal output
rlabel metal3 s 0 321104 800 321224 6 ch_data_out[72]
port 296 nsew signal output
rlabel metal3 s 0 320832 800 320952 6 ch_data_out[73]
port 297 nsew signal output
rlabel metal3 s 0 320560 800 320680 6 ch_data_out[74]
port 298 nsew signal output
rlabel metal3 s 0 320288 800 320408 6 ch_data_out[75]
port 299 nsew signal output
rlabel metal3 s 0 320016 800 320136 6 ch_data_out[76]
port 300 nsew signal output
rlabel metal3 s 59200 248616 60000 248736 6 ch_data_out[77]
port 301 nsew signal output
rlabel metal3 s 59200 248344 60000 248464 6 ch_data_out[78]
port 302 nsew signal output
rlabel metal3 s 59200 248072 60000 248192 6 ch_data_out[79]
port 303 nsew signal output
rlabel metal3 s 59200 1232 60000 1352 6 ch_data_out[7]
port 304 nsew signal output
rlabel metal3 s 59200 247800 60000 247920 6 ch_data_out[80]
port 305 nsew signal output
rlabel metal3 s 59200 247528 60000 247648 6 ch_data_out[81]
port 306 nsew signal output
rlabel metal3 s 59200 247256 60000 247376 6 ch_data_out[82]
port 307 nsew signal output
rlabel metal3 s 59200 246984 60000 247104 6 ch_data_out[83]
port 308 nsew signal output
rlabel metal3 s 59200 246712 60000 246832 6 ch_data_out[84]
port 309 nsew signal output
rlabel metal3 s 59200 246440 60000 246560 6 ch_data_out[85]
port 310 nsew signal output
rlabel metal3 s 59200 246168 60000 246288 6 ch_data_out[86]
port 311 nsew signal output
rlabel metal3 s 59200 245896 60000 246016 6 ch_data_out[87]
port 312 nsew signal output
rlabel metal3 s 59200 245624 60000 245744 6 ch_data_out[88]
port 313 nsew signal output
rlabel metal3 s 59200 245352 60000 245472 6 ch_data_out[89]
port 314 nsew signal output
rlabel metal3 s 59200 130840 60000 130960 6 ch_data_out[8]
port 315 nsew signal output
rlabel metal3 s 59200 245080 60000 245200 6 ch_data_out[90]
port 316 nsew signal output
rlabel metal3 s 59200 244808 60000 244928 6 ch_data_out[91]
port 317 nsew signal output
rlabel metal3 s 59200 244536 60000 244656 6 ch_data_out[92]
port 318 nsew signal output
rlabel metal3 s 59200 244264 60000 244384 6 ch_data_out[93]
port 319 nsew signal output
rlabel metal3 s 59200 243992 60000 244112 6 ch_data_out[94]
port 320 nsew signal output
rlabel metal3 s 59200 243720 60000 243840 6 ch_data_out[95]
port 321 nsew signal output
rlabel metal3 s 59200 243448 60000 243568 6 ch_data_out[96]
port 322 nsew signal output
rlabel metal3 s 59200 243176 60000 243296 6 ch_data_out[97]
port 323 nsew signal output
rlabel metal3 s 59200 242904 60000 243024 6 ch_data_out[98]
port 324 nsew signal output
rlabel metal3 s 59200 242632 60000 242752 6 ch_data_out[99]
port 325 nsew signal output
rlabel metal3 s 59200 130568 60000 130688 6 ch_data_out[9]
port 326 nsew signal output
rlabel metal2 s 13634 0 13690 800 6 clk_i
port 327 nsew signal input
rlabel metal2 s 38842 0 38898 800 6 m0_wbd_ack_o
port 328 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 m0_wbd_adr_i[0]
port 329 nsew signal input
rlabel metal2 s 24306 0 24362 800 6 m0_wbd_adr_i[10]
port 330 nsew signal input
rlabel metal2 s 24122 0 24178 800 6 m0_wbd_adr_i[11]
port 331 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 m0_wbd_adr_i[12]
port 332 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 m0_wbd_adr_i[13]
port 333 nsew signal input
rlabel metal2 s 23570 0 23626 800 6 m0_wbd_adr_i[14]
port 334 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 m0_wbd_adr_i[15]
port 335 nsew signal input
rlabel metal2 s 23202 0 23258 800 6 m0_wbd_adr_i[16]
port 336 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 m0_wbd_adr_i[17]
port 337 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 m0_wbd_adr_i[18]
port 338 nsew signal input
rlabel metal2 s 22650 0 22706 800 6 m0_wbd_adr_i[19]
port 339 nsew signal input
rlabel metal2 s 25962 0 26018 800 6 m0_wbd_adr_i[1]
port 340 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 m0_wbd_adr_i[20]
port 341 nsew signal input
rlabel metal2 s 22282 0 22338 800 6 m0_wbd_adr_i[21]
port 342 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 m0_wbd_adr_i[22]
port 343 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 m0_wbd_adr_i[23]
port 344 nsew signal input
rlabel metal2 s 21730 0 21786 800 6 m0_wbd_adr_i[24]
port 345 nsew signal input
rlabel metal2 s 21546 0 21602 800 6 m0_wbd_adr_i[25]
port 346 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 m0_wbd_adr_i[26]
port 347 nsew signal input
rlabel metal2 s 21178 0 21234 800 6 m0_wbd_adr_i[27]
port 348 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 m0_wbd_adr_i[28]
port 349 nsew signal input
rlabel metal2 s 20810 0 20866 800 6 m0_wbd_adr_i[29]
port 350 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 m0_wbd_adr_i[2]
port 351 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 m0_wbd_adr_i[30]
port 352 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 m0_wbd_adr_i[31]
port 353 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 m0_wbd_adr_i[3]
port 354 nsew signal input
rlabel metal2 s 25410 0 25466 800 6 m0_wbd_adr_i[4]
port 355 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 m0_wbd_adr_i[5]
port 356 nsew signal input
rlabel metal2 s 25042 0 25098 800 6 m0_wbd_adr_i[6]
port 357 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 m0_wbd_adr_i[7]
port 358 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 m0_wbd_adr_i[8]
port 359 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 m0_wbd_adr_i[9]
port 360 nsew signal input
rlabel metal2 s 39394 0 39450 800 6 m0_wbd_cyc_i
port 361 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 m0_wbd_dat_i[0]
port 362 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 m0_wbd_dat_i[10]
port 363 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 m0_wbd_dat_i[11]
port 364 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 m0_wbd_dat_i[12]
port 365 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 m0_wbd_dat_i[13]
port 366 nsew signal input
rlabel metal2 s 30194 0 30250 800 6 m0_wbd_dat_i[14]
port 367 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 m0_wbd_dat_i[15]
port 368 nsew signal input
rlabel metal2 s 29826 0 29882 800 6 m0_wbd_dat_i[16]
port 369 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 m0_wbd_dat_i[17]
port 370 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 m0_wbd_dat_i[18]
port 371 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 m0_wbd_dat_i[19]
port 372 nsew signal input
rlabel metal2 s 32586 0 32642 800 6 m0_wbd_dat_i[1]
port 373 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 m0_wbd_dat_i[20]
port 374 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 m0_wbd_dat_i[21]
port 375 nsew signal input
rlabel metal2 s 28722 0 28778 800 6 m0_wbd_dat_i[22]
port 376 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 m0_wbd_dat_i[23]
port 377 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 m0_wbd_dat_i[24]
port 378 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 m0_wbd_dat_i[25]
port 379 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 m0_wbd_dat_i[26]
port 380 nsew signal input
rlabel metal2 s 27802 0 27858 800 6 m0_wbd_dat_i[27]
port 381 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 m0_wbd_dat_i[28]
port 382 nsew signal input
rlabel metal2 s 27434 0 27490 800 6 m0_wbd_dat_i[29]
port 383 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 m0_wbd_dat_i[2]
port 384 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 m0_wbd_dat_i[30]
port 385 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 m0_wbd_dat_i[31]
port 386 nsew signal input
rlabel metal2 s 32218 0 32274 800 6 m0_wbd_dat_i[3]
port 387 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 m0_wbd_dat_i[4]
port 388 nsew signal input
rlabel metal2 s 31850 0 31906 800 6 m0_wbd_dat_i[5]
port 389 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 m0_wbd_dat_i[6]
port 390 nsew signal input
rlabel metal2 s 31482 0 31538 800 6 m0_wbd_dat_i[7]
port 391 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 m0_wbd_dat_i[8]
port 392 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 m0_wbd_dat_i[9]
port 393 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 m0_wbd_dat_o[0]
port 394 nsew signal output
rlabel metal2 s 36818 0 36874 800 6 m0_wbd_dat_o[10]
port 395 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 m0_wbd_dat_o[11]
port 396 nsew signal output
rlabel metal2 s 36450 0 36506 800 6 m0_wbd_dat_o[12]
port 397 nsew signal output
rlabel metal2 s 36266 0 36322 800 6 m0_wbd_dat_o[13]
port 398 nsew signal output
rlabel metal2 s 36082 0 36138 800 6 m0_wbd_dat_o[14]
port 399 nsew signal output
rlabel metal2 s 35898 0 35954 800 6 m0_wbd_dat_o[15]
port 400 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 m0_wbd_dat_o[16]
port 401 nsew signal output
rlabel metal2 s 35530 0 35586 800 6 m0_wbd_dat_o[17]
port 402 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 m0_wbd_dat_o[18]
port 403 nsew signal output
rlabel metal2 s 35162 0 35218 800 6 m0_wbd_dat_o[19]
port 404 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 m0_wbd_dat_o[1]
port 405 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 m0_wbd_dat_o[20]
port 406 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 m0_wbd_dat_o[21]
port 407 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 m0_wbd_dat_o[22]
port 408 nsew signal output
rlabel metal2 s 34426 0 34482 800 6 m0_wbd_dat_o[23]
port 409 nsew signal output
rlabel metal2 s 34242 0 34298 800 6 m0_wbd_dat_o[24]
port 410 nsew signal output
rlabel metal2 s 34058 0 34114 800 6 m0_wbd_dat_o[25]
port 411 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 m0_wbd_dat_o[26]
port 412 nsew signal output
rlabel metal2 s 33690 0 33746 800 6 m0_wbd_dat_o[27]
port 413 nsew signal output
rlabel metal2 s 33506 0 33562 800 6 m0_wbd_dat_o[28]
port 414 nsew signal output
rlabel metal2 s 33322 0 33378 800 6 m0_wbd_dat_o[29]
port 415 nsew signal output
rlabel metal2 s 38290 0 38346 800 6 m0_wbd_dat_o[2]
port 416 nsew signal output
rlabel metal2 s 33138 0 33194 800 6 m0_wbd_dat_o[30]
port 417 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 m0_wbd_dat_o[31]
port 418 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 m0_wbd_dat_o[3]
port 419 nsew signal output
rlabel metal2 s 37922 0 37978 800 6 m0_wbd_dat_o[4]
port 420 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 m0_wbd_dat_o[5]
port 421 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 m0_wbd_dat_o[6]
port 422 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 m0_wbd_dat_o[7]
port 423 nsew signal output
rlabel metal2 s 37186 0 37242 800 6 m0_wbd_dat_o[8]
port 424 nsew signal output
rlabel metal2 s 37002 0 37058 800 6 m0_wbd_dat_o[9]
port 425 nsew signal output
rlabel metal2 s 39210 0 39266 800 6 m0_wbd_err_o
port 426 nsew signal output
rlabel metal2 s 39026 0 39082 800 6 m0_wbd_lack_o
port 427 nsew signal output
rlabel metal2 s 26882 0 26938 800 6 m0_wbd_sel_i[0]
port 428 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 m0_wbd_sel_i[1]
port 429 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 m0_wbd_sel_i[2]
port 430 nsew signal input
rlabel metal2 s 26330 0 26386 800 6 m0_wbd_sel_i[3]
port 431 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 m0_wbd_stb_i
port 432 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 m0_wbd_we_i
port 433 nsew signal input
rlabel metal3 s 0 49512 800 49632 6 m1_wbd_ack_o
port 434 nsew signal output
rlabel metal3 s 0 29384 800 29504 6 m1_wbd_adr_i[0]
port 435 nsew signal input
rlabel metal3 s 0 26664 800 26784 6 m1_wbd_adr_i[10]
port 436 nsew signal input
rlabel metal3 s 0 26392 800 26512 6 m1_wbd_adr_i[11]
port 437 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 m1_wbd_adr_i[12]
port 438 nsew signal input
rlabel metal3 s 0 25848 800 25968 6 m1_wbd_adr_i[13]
port 439 nsew signal input
rlabel metal3 s 0 25576 800 25696 6 m1_wbd_adr_i[14]
port 440 nsew signal input
rlabel metal3 s 0 25304 800 25424 6 m1_wbd_adr_i[15]
port 441 nsew signal input
rlabel metal3 s 0 25032 800 25152 6 m1_wbd_adr_i[16]
port 442 nsew signal input
rlabel metal3 s 0 24760 800 24880 6 m1_wbd_adr_i[17]
port 443 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 m1_wbd_adr_i[18]
port 444 nsew signal input
rlabel metal3 s 0 24216 800 24336 6 m1_wbd_adr_i[19]
port 445 nsew signal input
rlabel metal3 s 0 29112 800 29232 6 m1_wbd_adr_i[1]
port 446 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 m1_wbd_adr_i[20]
port 447 nsew signal input
rlabel metal3 s 0 23672 800 23792 6 m1_wbd_adr_i[21]
port 448 nsew signal input
rlabel metal3 s 0 23400 800 23520 6 m1_wbd_adr_i[22]
port 449 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 m1_wbd_adr_i[23]
port 450 nsew signal input
rlabel metal3 s 0 22856 800 22976 6 m1_wbd_adr_i[24]
port 451 nsew signal input
rlabel metal3 s 0 22584 800 22704 6 m1_wbd_adr_i[25]
port 452 nsew signal input
rlabel metal3 s 0 22312 800 22432 6 m1_wbd_adr_i[26]
port 453 nsew signal input
rlabel metal3 s 0 22040 800 22160 6 m1_wbd_adr_i[27]
port 454 nsew signal input
rlabel metal3 s 0 21768 800 21888 6 m1_wbd_adr_i[28]
port 455 nsew signal input
rlabel metal3 s 0 21496 800 21616 6 m1_wbd_adr_i[29]
port 456 nsew signal input
rlabel metal3 s 0 28840 800 28960 6 m1_wbd_adr_i[2]
port 457 nsew signal input
rlabel metal3 s 0 21224 800 21344 6 m1_wbd_adr_i[30]
port 458 nsew signal input
rlabel metal3 s 0 20952 800 21072 6 m1_wbd_adr_i[31]
port 459 nsew signal input
rlabel metal3 s 0 28568 800 28688 6 m1_wbd_adr_i[3]
port 460 nsew signal input
rlabel metal3 s 0 28296 800 28416 6 m1_wbd_adr_i[4]
port 461 nsew signal input
rlabel metal3 s 0 28024 800 28144 6 m1_wbd_adr_i[5]
port 462 nsew signal input
rlabel metal3 s 0 27752 800 27872 6 m1_wbd_adr_i[6]
port 463 nsew signal input
rlabel metal3 s 0 27480 800 27600 6 m1_wbd_adr_i[7]
port 464 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 m1_wbd_adr_i[8]
port 465 nsew signal input
rlabel metal3 s 0 26936 800 27056 6 m1_wbd_adr_i[9]
port 466 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 m1_wbd_bl_i[0]
port 467 nsew signal input
rlabel metal3 s 0 31016 800 31136 6 m1_wbd_bl_i[1]
port 468 nsew signal input
rlabel metal3 s 0 30744 800 30864 6 m1_wbd_bl_i[2]
port 469 nsew signal input
rlabel metal3 s 0 31560 800 31680 6 m1_wbd_bry_i
port 470 nsew signal input
rlabel metal3 s 0 20408 800 20528 6 m1_wbd_cyc_i
port 471 nsew signal input
rlabel metal3 s 0 40264 800 40384 6 m1_wbd_dat_i[0]
port 472 nsew signal input
rlabel metal3 s 0 37544 800 37664 6 m1_wbd_dat_i[10]
port 473 nsew signal input
rlabel metal3 s 0 37272 800 37392 6 m1_wbd_dat_i[11]
port 474 nsew signal input
rlabel metal3 s 0 37000 800 37120 6 m1_wbd_dat_i[12]
port 475 nsew signal input
rlabel metal3 s 0 36728 800 36848 6 m1_wbd_dat_i[13]
port 476 nsew signal input
rlabel metal3 s 0 36456 800 36576 6 m1_wbd_dat_i[14]
port 477 nsew signal input
rlabel metal3 s 0 36184 800 36304 6 m1_wbd_dat_i[15]
port 478 nsew signal input
rlabel metal3 s 0 35912 800 36032 6 m1_wbd_dat_i[16]
port 479 nsew signal input
rlabel metal3 s 0 35640 800 35760 6 m1_wbd_dat_i[17]
port 480 nsew signal input
rlabel metal3 s 0 35368 800 35488 6 m1_wbd_dat_i[18]
port 481 nsew signal input
rlabel metal3 s 0 35096 800 35216 6 m1_wbd_dat_i[19]
port 482 nsew signal input
rlabel metal3 s 0 39992 800 40112 6 m1_wbd_dat_i[1]
port 483 nsew signal input
rlabel metal3 s 0 34824 800 34944 6 m1_wbd_dat_i[20]
port 484 nsew signal input
rlabel metal3 s 0 34552 800 34672 6 m1_wbd_dat_i[21]
port 485 nsew signal input
rlabel metal3 s 0 34280 800 34400 6 m1_wbd_dat_i[22]
port 486 nsew signal input
rlabel metal3 s 0 34008 800 34128 6 m1_wbd_dat_i[23]
port 487 nsew signal input
rlabel metal3 s 0 33736 800 33856 6 m1_wbd_dat_i[24]
port 488 nsew signal input
rlabel metal3 s 0 33464 800 33584 6 m1_wbd_dat_i[25]
port 489 nsew signal input
rlabel metal3 s 0 33192 800 33312 6 m1_wbd_dat_i[26]
port 490 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 m1_wbd_dat_i[27]
port 491 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 m1_wbd_dat_i[28]
port 492 nsew signal input
rlabel metal3 s 0 32376 800 32496 6 m1_wbd_dat_i[29]
port 493 nsew signal input
rlabel metal3 s 0 39720 800 39840 6 m1_wbd_dat_i[2]
port 494 nsew signal input
rlabel metal3 s 0 32104 800 32224 6 m1_wbd_dat_i[30]
port 495 nsew signal input
rlabel metal3 s 0 31832 800 31952 6 m1_wbd_dat_i[31]
port 496 nsew signal input
rlabel metal3 s 0 39448 800 39568 6 m1_wbd_dat_i[3]
port 497 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 m1_wbd_dat_i[4]
port 498 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 m1_wbd_dat_i[5]
port 499 nsew signal input
rlabel metal3 s 0 38632 800 38752 6 m1_wbd_dat_i[6]
port 500 nsew signal input
rlabel metal3 s 0 38360 800 38480 6 m1_wbd_dat_i[7]
port 501 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 m1_wbd_dat_i[8]
port 502 nsew signal input
rlabel metal3 s 0 37816 800 37936 6 m1_wbd_dat_i[9]
port 503 nsew signal input
rlabel metal3 s 0 48968 800 49088 6 m1_wbd_dat_o[0]
port 504 nsew signal output
rlabel metal3 s 0 46248 800 46368 6 m1_wbd_dat_o[10]
port 505 nsew signal output
rlabel metal3 s 0 45976 800 46096 6 m1_wbd_dat_o[11]
port 506 nsew signal output
rlabel metal3 s 0 45704 800 45824 6 m1_wbd_dat_o[12]
port 507 nsew signal output
rlabel metal3 s 0 45432 800 45552 6 m1_wbd_dat_o[13]
port 508 nsew signal output
rlabel metal3 s 0 45160 800 45280 6 m1_wbd_dat_o[14]
port 509 nsew signal output
rlabel metal3 s 0 44888 800 45008 6 m1_wbd_dat_o[15]
port 510 nsew signal output
rlabel metal3 s 0 44616 800 44736 6 m1_wbd_dat_o[16]
port 511 nsew signal output
rlabel metal3 s 0 44344 800 44464 6 m1_wbd_dat_o[17]
port 512 nsew signal output
rlabel metal3 s 0 44072 800 44192 6 m1_wbd_dat_o[18]
port 513 nsew signal output
rlabel metal3 s 0 43800 800 43920 6 m1_wbd_dat_o[19]
port 514 nsew signal output
rlabel metal3 s 0 48696 800 48816 6 m1_wbd_dat_o[1]
port 515 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 m1_wbd_dat_o[20]
port 516 nsew signal output
rlabel metal3 s 0 43256 800 43376 6 m1_wbd_dat_o[21]
port 517 nsew signal output
rlabel metal3 s 0 42984 800 43104 6 m1_wbd_dat_o[22]
port 518 nsew signal output
rlabel metal3 s 0 42712 800 42832 6 m1_wbd_dat_o[23]
port 519 nsew signal output
rlabel metal3 s 0 42440 800 42560 6 m1_wbd_dat_o[24]
port 520 nsew signal output
rlabel metal3 s 0 42168 800 42288 6 m1_wbd_dat_o[25]
port 521 nsew signal output
rlabel metal3 s 0 41896 800 42016 6 m1_wbd_dat_o[26]
port 522 nsew signal output
rlabel metal3 s 0 41624 800 41744 6 m1_wbd_dat_o[27]
port 523 nsew signal output
rlabel metal3 s 0 41352 800 41472 6 m1_wbd_dat_o[28]
port 524 nsew signal output
rlabel metal3 s 0 41080 800 41200 6 m1_wbd_dat_o[29]
port 525 nsew signal output
rlabel metal3 s 0 48424 800 48544 6 m1_wbd_dat_o[2]
port 526 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 m1_wbd_dat_o[30]
port 527 nsew signal output
rlabel metal3 s 0 40536 800 40656 6 m1_wbd_dat_o[31]
port 528 nsew signal output
rlabel metal3 s 0 48152 800 48272 6 m1_wbd_dat_o[3]
port 529 nsew signal output
rlabel metal3 s 0 47880 800 48000 6 m1_wbd_dat_o[4]
port 530 nsew signal output
rlabel metal3 s 0 47608 800 47728 6 m1_wbd_dat_o[5]
port 531 nsew signal output
rlabel metal3 s 0 47336 800 47456 6 m1_wbd_dat_o[6]
port 532 nsew signal output
rlabel metal3 s 0 47064 800 47184 6 m1_wbd_dat_o[7]
port 533 nsew signal output
rlabel metal3 s 0 46792 800 46912 6 m1_wbd_dat_o[8]
port 534 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 m1_wbd_dat_o[9]
port 535 nsew signal output
rlabel metal3 s 0 49784 800 49904 6 m1_wbd_err_o
port 536 nsew signal output
rlabel metal3 s 0 49240 800 49360 6 m1_wbd_lack_o
port 537 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 m1_wbd_sel_i[0]
port 538 nsew signal input
rlabel metal3 s 0 30200 800 30320 6 m1_wbd_sel_i[1]
port 539 nsew signal input
rlabel metal3 s 0 29928 800 30048 6 m1_wbd_sel_i[2]
port 540 nsew signal input
rlabel metal3 s 0 29656 800 29776 6 m1_wbd_sel_i[3]
port 541 nsew signal input
rlabel metal3 s 0 20136 800 20256 6 m1_wbd_stb_i
port 542 nsew signal input
rlabel metal3 s 0 20680 800 20800 6 m1_wbd_we_i
port 543 nsew signal input
rlabel metal3 s 0 91128 800 91248 6 m2_wbd_ack_o
port 544 nsew signal output
rlabel metal3 s 0 69368 800 69488 6 m2_wbd_adr_i[0]
port 545 nsew signal input
rlabel metal3 s 0 66648 800 66768 6 m2_wbd_adr_i[10]
port 546 nsew signal input
rlabel metal3 s 0 66376 800 66496 6 m2_wbd_adr_i[11]
port 547 nsew signal input
rlabel metal3 s 0 66104 800 66224 6 m2_wbd_adr_i[12]
port 548 nsew signal input
rlabel metal3 s 0 65832 800 65952 6 m2_wbd_adr_i[13]
port 549 nsew signal input
rlabel metal3 s 0 65560 800 65680 6 m2_wbd_adr_i[14]
port 550 nsew signal input
rlabel metal3 s 0 65288 800 65408 6 m2_wbd_adr_i[15]
port 551 nsew signal input
rlabel metal3 s 0 65016 800 65136 6 m2_wbd_adr_i[16]
port 552 nsew signal input
rlabel metal3 s 0 64744 800 64864 6 m2_wbd_adr_i[17]
port 553 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 m2_wbd_adr_i[18]
port 554 nsew signal input
rlabel metal3 s 0 64200 800 64320 6 m2_wbd_adr_i[19]
port 555 nsew signal input
rlabel metal3 s 0 69096 800 69216 6 m2_wbd_adr_i[1]
port 556 nsew signal input
rlabel metal3 s 0 63928 800 64048 6 m2_wbd_adr_i[20]
port 557 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 m2_wbd_adr_i[21]
port 558 nsew signal input
rlabel metal3 s 0 63384 800 63504 6 m2_wbd_adr_i[22]
port 559 nsew signal input
rlabel metal3 s 0 63112 800 63232 6 m2_wbd_adr_i[23]
port 560 nsew signal input
rlabel metal3 s 0 62840 800 62960 6 m2_wbd_adr_i[24]
port 561 nsew signal input
rlabel metal3 s 0 62568 800 62688 6 m2_wbd_adr_i[25]
port 562 nsew signal input
rlabel metal3 s 0 62296 800 62416 6 m2_wbd_adr_i[26]
port 563 nsew signal input
rlabel metal3 s 0 62024 800 62144 6 m2_wbd_adr_i[27]
port 564 nsew signal input
rlabel metal3 s 0 61752 800 61872 6 m2_wbd_adr_i[28]
port 565 nsew signal input
rlabel metal3 s 0 61480 800 61600 6 m2_wbd_adr_i[29]
port 566 nsew signal input
rlabel metal3 s 0 68824 800 68944 6 m2_wbd_adr_i[2]
port 567 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 m2_wbd_adr_i[30]
port 568 nsew signal input
rlabel metal3 s 0 60936 800 61056 6 m2_wbd_adr_i[31]
port 569 nsew signal input
rlabel metal3 s 0 68552 800 68672 6 m2_wbd_adr_i[3]
port 570 nsew signal input
rlabel metal3 s 0 68280 800 68400 6 m2_wbd_adr_i[4]
port 571 nsew signal input
rlabel metal3 s 0 68008 800 68128 6 m2_wbd_adr_i[5]
port 572 nsew signal input
rlabel metal3 s 0 67736 800 67856 6 m2_wbd_adr_i[6]
port 573 nsew signal input
rlabel metal3 s 0 67464 800 67584 6 m2_wbd_adr_i[7]
port 574 nsew signal input
rlabel metal3 s 0 67192 800 67312 6 m2_wbd_adr_i[8]
port 575 nsew signal input
rlabel metal3 s 0 66920 800 67040 6 m2_wbd_adr_i[9]
port 576 nsew signal input
rlabel metal3 s 0 73176 800 73296 6 m2_wbd_bl_i[0]
port 577 nsew signal input
rlabel metal3 s 0 72904 800 73024 6 m2_wbd_bl_i[1]
port 578 nsew signal input
rlabel metal3 s 0 72632 800 72752 6 m2_wbd_bl_i[2]
port 579 nsew signal input
rlabel metal3 s 0 72360 800 72480 6 m2_wbd_bl_i[3]
port 580 nsew signal input
rlabel metal3 s 0 72088 800 72208 6 m2_wbd_bl_i[4]
port 581 nsew signal input
rlabel metal3 s 0 71816 800 71936 6 m2_wbd_bl_i[5]
port 582 nsew signal input
rlabel metal3 s 0 71544 800 71664 6 m2_wbd_bl_i[6]
port 583 nsew signal input
rlabel metal3 s 0 71272 800 71392 6 m2_wbd_bl_i[7]
port 584 nsew signal input
rlabel metal3 s 0 71000 800 71120 6 m2_wbd_bl_i[8]
port 585 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 m2_wbd_bl_i[9]
port 586 nsew signal input
rlabel metal3 s 0 73448 800 73568 6 m2_wbd_bry_i
port 587 nsew signal input
rlabel metal3 s 0 60392 800 60512 6 m2_wbd_cyc_i
port 588 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 m2_wbd_dat_i[0]
port 589 nsew signal input
rlabel metal3 s 0 79432 800 79552 6 m2_wbd_dat_i[10]
port 590 nsew signal input
rlabel metal3 s 0 79160 800 79280 6 m2_wbd_dat_i[11]
port 591 nsew signal input
rlabel metal3 s 0 78888 800 79008 6 m2_wbd_dat_i[12]
port 592 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 m2_wbd_dat_i[13]
port 593 nsew signal input
rlabel metal3 s 0 78344 800 78464 6 m2_wbd_dat_i[14]
port 594 nsew signal input
rlabel metal3 s 0 78072 800 78192 6 m2_wbd_dat_i[15]
port 595 nsew signal input
rlabel metal3 s 0 77800 800 77920 6 m2_wbd_dat_i[16]
port 596 nsew signal input
rlabel metal3 s 0 77528 800 77648 6 m2_wbd_dat_i[17]
port 597 nsew signal input
rlabel metal3 s 0 77256 800 77376 6 m2_wbd_dat_i[18]
port 598 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 m2_wbd_dat_i[19]
port 599 nsew signal input
rlabel metal3 s 0 81880 800 82000 6 m2_wbd_dat_i[1]
port 600 nsew signal input
rlabel metal3 s 0 76712 800 76832 6 m2_wbd_dat_i[20]
port 601 nsew signal input
rlabel metal3 s 0 76440 800 76560 6 m2_wbd_dat_i[21]
port 602 nsew signal input
rlabel metal3 s 0 76168 800 76288 6 m2_wbd_dat_i[22]
port 603 nsew signal input
rlabel metal3 s 0 75896 800 76016 6 m2_wbd_dat_i[23]
port 604 nsew signal input
rlabel metal3 s 0 75624 800 75744 6 m2_wbd_dat_i[24]
port 605 nsew signal input
rlabel metal3 s 0 75352 800 75472 6 m2_wbd_dat_i[25]
port 606 nsew signal input
rlabel metal3 s 0 75080 800 75200 6 m2_wbd_dat_i[26]
port 607 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 m2_wbd_dat_i[27]
port 608 nsew signal input
rlabel metal3 s 0 74536 800 74656 6 m2_wbd_dat_i[28]
port 609 nsew signal input
rlabel metal3 s 0 74264 800 74384 6 m2_wbd_dat_i[29]
port 610 nsew signal input
rlabel metal3 s 0 81608 800 81728 6 m2_wbd_dat_i[2]
port 611 nsew signal input
rlabel metal3 s 0 73992 800 74112 6 m2_wbd_dat_i[30]
port 612 nsew signal input
rlabel metal3 s 0 73720 800 73840 6 m2_wbd_dat_i[31]
port 613 nsew signal input
rlabel metal3 s 0 81336 800 81456 6 m2_wbd_dat_i[3]
port 614 nsew signal input
rlabel metal3 s 0 81064 800 81184 6 m2_wbd_dat_i[4]
port 615 nsew signal input
rlabel metal3 s 0 80792 800 80912 6 m2_wbd_dat_i[5]
port 616 nsew signal input
rlabel metal3 s 0 80520 800 80640 6 m2_wbd_dat_i[6]
port 617 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 m2_wbd_dat_i[7]
port 618 nsew signal input
rlabel metal3 s 0 79976 800 80096 6 m2_wbd_dat_i[8]
port 619 nsew signal input
rlabel metal3 s 0 79704 800 79824 6 m2_wbd_dat_i[9]
port 620 nsew signal input
rlabel metal3 s 0 90856 800 90976 6 m2_wbd_dat_o[0]
port 621 nsew signal output
rlabel metal3 s 0 88136 800 88256 6 m2_wbd_dat_o[10]
port 622 nsew signal output
rlabel metal3 s 0 87864 800 87984 6 m2_wbd_dat_o[11]
port 623 nsew signal output
rlabel metal3 s 0 87592 800 87712 6 m2_wbd_dat_o[12]
port 624 nsew signal output
rlabel metal3 s 0 87320 800 87440 6 m2_wbd_dat_o[13]
port 625 nsew signal output
rlabel metal3 s 0 87048 800 87168 6 m2_wbd_dat_o[14]
port 626 nsew signal output
rlabel metal3 s 0 86776 800 86896 6 m2_wbd_dat_o[15]
port 627 nsew signal output
rlabel metal3 s 0 86504 800 86624 6 m2_wbd_dat_o[16]
port 628 nsew signal output
rlabel metal3 s 0 86232 800 86352 6 m2_wbd_dat_o[17]
port 629 nsew signal output
rlabel metal3 s 0 85960 800 86080 6 m2_wbd_dat_o[18]
port 630 nsew signal output
rlabel metal3 s 0 85688 800 85808 6 m2_wbd_dat_o[19]
port 631 nsew signal output
rlabel metal3 s 0 90584 800 90704 6 m2_wbd_dat_o[1]
port 632 nsew signal output
rlabel metal3 s 0 85416 800 85536 6 m2_wbd_dat_o[20]
port 633 nsew signal output
rlabel metal3 s 0 85144 800 85264 6 m2_wbd_dat_o[21]
port 634 nsew signal output
rlabel metal3 s 0 84872 800 84992 6 m2_wbd_dat_o[22]
port 635 nsew signal output
rlabel metal3 s 0 84600 800 84720 6 m2_wbd_dat_o[23]
port 636 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 m2_wbd_dat_o[24]
port 637 nsew signal output
rlabel metal3 s 0 84056 800 84176 6 m2_wbd_dat_o[25]
port 638 nsew signal output
rlabel metal3 s 0 83784 800 83904 6 m2_wbd_dat_o[26]
port 639 nsew signal output
rlabel metal3 s 0 83512 800 83632 6 m2_wbd_dat_o[27]
port 640 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 m2_wbd_dat_o[28]
port 641 nsew signal output
rlabel metal3 s 0 82968 800 83088 6 m2_wbd_dat_o[29]
port 642 nsew signal output
rlabel metal3 s 0 90312 800 90432 6 m2_wbd_dat_o[2]
port 643 nsew signal output
rlabel metal3 s 0 82696 800 82816 6 m2_wbd_dat_o[30]
port 644 nsew signal output
rlabel metal3 s 0 82424 800 82544 6 m2_wbd_dat_o[31]
port 645 nsew signal output
rlabel metal3 s 0 90040 800 90160 6 m2_wbd_dat_o[3]
port 646 nsew signal output
rlabel metal3 s 0 89768 800 89888 6 m2_wbd_dat_o[4]
port 647 nsew signal output
rlabel metal3 s 0 89496 800 89616 6 m2_wbd_dat_o[5]
port 648 nsew signal output
rlabel metal3 s 0 89224 800 89344 6 m2_wbd_dat_o[6]
port 649 nsew signal output
rlabel metal3 s 0 88952 800 89072 6 m2_wbd_dat_o[7]
port 650 nsew signal output
rlabel metal3 s 0 88680 800 88800 6 m2_wbd_dat_o[8]
port 651 nsew signal output
rlabel metal3 s 0 88408 800 88528 6 m2_wbd_dat_o[9]
port 652 nsew signal output
rlabel metal3 s 0 91672 800 91792 6 m2_wbd_err_o
port 653 nsew signal output
rlabel metal3 s 0 91400 800 91520 6 m2_wbd_lack_o
port 654 nsew signal output
rlabel metal3 s 0 70456 800 70576 6 m2_wbd_sel_i[0]
port 655 nsew signal input
rlabel metal3 s 0 70184 800 70304 6 m2_wbd_sel_i[1]
port 656 nsew signal input
rlabel metal3 s 0 69912 800 70032 6 m2_wbd_sel_i[2]
port 657 nsew signal input
rlabel metal3 s 0 69640 800 69760 6 m2_wbd_sel_i[3]
port 658 nsew signal input
rlabel metal3 s 0 60120 800 60240 6 m2_wbd_stb_i
port 659 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 m2_wbd_we_i
port 660 nsew signal input
rlabel metal3 s 0 122408 800 122528 6 m3_wbd_ack_o
port 661 nsew signal output
rlabel metal3 s 0 109352 800 109472 6 m3_wbd_adr_i[0]
port 662 nsew signal input
rlabel metal3 s 0 106632 800 106752 6 m3_wbd_adr_i[10]
port 663 nsew signal input
rlabel metal3 s 0 106360 800 106480 6 m3_wbd_adr_i[11]
port 664 nsew signal input
rlabel metal3 s 0 106088 800 106208 6 m3_wbd_adr_i[12]
port 665 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 m3_wbd_adr_i[13]
port 666 nsew signal input
rlabel metal3 s 0 105544 800 105664 6 m3_wbd_adr_i[14]
port 667 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 m3_wbd_adr_i[15]
port 668 nsew signal input
rlabel metal3 s 0 105000 800 105120 6 m3_wbd_adr_i[16]
port 669 nsew signal input
rlabel metal3 s 0 104728 800 104848 6 m3_wbd_adr_i[17]
port 670 nsew signal input
rlabel metal3 s 0 104456 800 104576 6 m3_wbd_adr_i[18]
port 671 nsew signal input
rlabel metal3 s 0 104184 800 104304 6 m3_wbd_adr_i[19]
port 672 nsew signal input
rlabel metal3 s 0 109080 800 109200 6 m3_wbd_adr_i[1]
port 673 nsew signal input
rlabel metal3 s 0 103912 800 104032 6 m3_wbd_adr_i[20]
port 674 nsew signal input
rlabel metal3 s 0 103640 800 103760 6 m3_wbd_adr_i[21]
port 675 nsew signal input
rlabel metal3 s 0 103368 800 103488 6 m3_wbd_adr_i[22]
port 676 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 m3_wbd_adr_i[23]
port 677 nsew signal input
rlabel metal3 s 0 102824 800 102944 6 m3_wbd_adr_i[24]
port 678 nsew signal input
rlabel metal3 s 0 102552 800 102672 6 m3_wbd_adr_i[25]
port 679 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 m3_wbd_adr_i[26]
port 680 nsew signal input
rlabel metal3 s 0 102008 800 102128 6 m3_wbd_adr_i[27]
port 681 nsew signal input
rlabel metal3 s 0 101736 800 101856 6 m3_wbd_adr_i[28]
port 682 nsew signal input
rlabel metal3 s 0 101464 800 101584 6 m3_wbd_adr_i[29]
port 683 nsew signal input
rlabel metal3 s 0 108808 800 108928 6 m3_wbd_adr_i[2]
port 684 nsew signal input
rlabel metal3 s 0 101192 800 101312 6 m3_wbd_adr_i[30]
port 685 nsew signal input
rlabel metal3 s 0 100920 800 101040 6 m3_wbd_adr_i[31]
port 686 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 m3_wbd_adr_i[3]
port 687 nsew signal input
rlabel metal3 s 0 108264 800 108384 6 m3_wbd_adr_i[4]
port 688 nsew signal input
rlabel metal3 s 0 107992 800 108112 6 m3_wbd_adr_i[5]
port 689 nsew signal input
rlabel metal3 s 0 107720 800 107840 6 m3_wbd_adr_i[6]
port 690 nsew signal input
rlabel metal3 s 0 107448 800 107568 6 m3_wbd_adr_i[7]
port 691 nsew signal input
rlabel metal3 s 0 107176 800 107296 6 m3_wbd_adr_i[8]
port 692 nsew signal input
rlabel metal3 s 0 106904 800 107024 6 m3_wbd_adr_i[9]
port 693 nsew signal input
rlabel metal3 s 0 113160 800 113280 6 m3_wbd_bl_i[0]
port 694 nsew signal input
rlabel metal3 s 0 112888 800 113008 6 m3_wbd_bl_i[1]
port 695 nsew signal input
rlabel metal3 s 0 112616 800 112736 6 m3_wbd_bl_i[2]
port 696 nsew signal input
rlabel metal3 s 0 112344 800 112464 6 m3_wbd_bl_i[3]
port 697 nsew signal input
rlabel metal3 s 0 112072 800 112192 6 m3_wbd_bl_i[4]
port 698 nsew signal input
rlabel metal3 s 0 111800 800 111920 6 m3_wbd_bl_i[5]
port 699 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 m3_wbd_bl_i[6]
port 700 nsew signal input
rlabel metal3 s 0 111256 800 111376 6 m3_wbd_bl_i[7]
port 701 nsew signal input
rlabel metal3 s 0 110984 800 111104 6 m3_wbd_bl_i[8]
port 702 nsew signal input
rlabel metal3 s 0 110712 800 110832 6 m3_wbd_bl_i[9]
port 703 nsew signal input
rlabel metal3 s 0 113432 800 113552 6 m3_wbd_bry_i
port 704 nsew signal input
rlabel metal3 s 0 100376 800 100496 6 m3_wbd_cyc_i
port 705 nsew signal input
rlabel metal3 s 0 122136 800 122256 6 m3_wbd_dat_o[0]
port 706 nsew signal output
rlabel metal3 s 0 119416 800 119536 6 m3_wbd_dat_o[10]
port 707 nsew signal output
rlabel metal3 s 0 119144 800 119264 6 m3_wbd_dat_o[11]
port 708 nsew signal output
rlabel metal3 s 0 118872 800 118992 6 m3_wbd_dat_o[12]
port 709 nsew signal output
rlabel metal3 s 0 118600 800 118720 6 m3_wbd_dat_o[13]
port 710 nsew signal output
rlabel metal3 s 0 118328 800 118448 6 m3_wbd_dat_o[14]
port 711 nsew signal output
rlabel metal3 s 0 118056 800 118176 6 m3_wbd_dat_o[15]
port 712 nsew signal output
rlabel metal3 s 0 117784 800 117904 6 m3_wbd_dat_o[16]
port 713 nsew signal output
rlabel metal3 s 0 117512 800 117632 6 m3_wbd_dat_o[17]
port 714 nsew signal output
rlabel metal3 s 0 117240 800 117360 6 m3_wbd_dat_o[18]
port 715 nsew signal output
rlabel metal3 s 0 116968 800 117088 6 m3_wbd_dat_o[19]
port 716 nsew signal output
rlabel metal3 s 0 121864 800 121984 6 m3_wbd_dat_o[1]
port 717 nsew signal output
rlabel metal3 s 0 116696 800 116816 6 m3_wbd_dat_o[20]
port 718 nsew signal output
rlabel metal3 s 0 116424 800 116544 6 m3_wbd_dat_o[21]
port 719 nsew signal output
rlabel metal3 s 0 116152 800 116272 6 m3_wbd_dat_o[22]
port 720 nsew signal output
rlabel metal3 s 0 115880 800 116000 6 m3_wbd_dat_o[23]
port 721 nsew signal output
rlabel metal3 s 0 115608 800 115728 6 m3_wbd_dat_o[24]
port 722 nsew signal output
rlabel metal3 s 0 115336 800 115456 6 m3_wbd_dat_o[25]
port 723 nsew signal output
rlabel metal3 s 0 115064 800 115184 6 m3_wbd_dat_o[26]
port 724 nsew signal output
rlabel metal3 s 0 114792 800 114912 6 m3_wbd_dat_o[27]
port 725 nsew signal output
rlabel metal3 s 0 114520 800 114640 6 m3_wbd_dat_o[28]
port 726 nsew signal output
rlabel metal3 s 0 114248 800 114368 6 m3_wbd_dat_o[29]
port 727 nsew signal output
rlabel metal3 s 0 121592 800 121712 6 m3_wbd_dat_o[2]
port 728 nsew signal output
rlabel metal3 s 0 113976 800 114096 6 m3_wbd_dat_o[30]
port 729 nsew signal output
rlabel metal3 s 0 113704 800 113824 6 m3_wbd_dat_o[31]
port 730 nsew signal output
rlabel metal3 s 0 121320 800 121440 6 m3_wbd_dat_o[3]
port 731 nsew signal output
rlabel metal3 s 0 121048 800 121168 6 m3_wbd_dat_o[4]
port 732 nsew signal output
rlabel metal3 s 0 120776 800 120896 6 m3_wbd_dat_o[5]
port 733 nsew signal output
rlabel metal3 s 0 120504 800 120624 6 m3_wbd_dat_o[6]
port 734 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 m3_wbd_dat_o[7]
port 735 nsew signal output
rlabel metal3 s 0 119960 800 120080 6 m3_wbd_dat_o[8]
port 736 nsew signal output
rlabel metal3 s 0 119688 800 119808 6 m3_wbd_dat_o[9]
port 737 nsew signal output
rlabel metal3 s 0 122952 800 123072 6 m3_wbd_err_o
port 738 nsew signal output
rlabel metal3 s 0 122680 800 122800 6 m3_wbd_lack_o
port 739 nsew signal output
rlabel metal3 s 0 110440 800 110560 6 m3_wbd_sel_i[0]
port 740 nsew signal input
rlabel metal3 s 0 110168 800 110288 6 m3_wbd_sel_i[1]
port 741 nsew signal input
rlabel metal3 s 0 109896 800 110016 6 m3_wbd_sel_i[2]
port 742 nsew signal input
rlabel metal3 s 0 109624 800 109744 6 m3_wbd_sel_i[3]
port 743 nsew signal input
rlabel metal3 s 0 100104 800 100224 6 m3_wbd_stb_i
port 744 nsew signal input
rlabel metal3 s 0 100648 800 100768 6 m3_wbd_we_i
port 745 nsew signal input
rlabel metal2 s 13082 0 13138 800 6 mclk_raw
port 746 nsew signal input
rlabel metal3 s 59200 350072 60000 350192 6 peri_wbclk
port 747 nsew signal output
rlabel metal3 s 0 11160 800 11280 6 riscv_wbclk
port 748 nsew signal output
rlabel metal2 s 4066 0 4122 800 6 rst_n
port 749 nsew signal input
rlabel metal3 s 59200 10344 60000 10464 6 s0_idle
port 750 nsew signal input
rlabel metal3 s 59200 10072 60000 10192 6 s0_mclk
port 751 nsew signal output
rlabel metal3 s 59200 41352 60000 41472 6 s0_wbd_ack_i
port 752 nsew signal input
rlabel metal3 s 59200 19592 60000 19712 6 s0_wbd_adr_o[0]
port 753 nsew signal output
rlabel metal3 s 59200 16872 60000 16992 6 s0_wbd_adr_o[10]
port 754 nsew signal output
rlabel metal3 s 59200 16600 60000 16720 6 s0_wbd_adr_o[11]
port 755 nsew signal output
rlabel metal3 s 59200 16328 60000 16448 6 s0_wbd_adr_o[12]
port 756 nsew signal output
rlabel metal3 s 59200 16056 60000 16176 6 s0_wbd_adr_o[13]
port 757 nsew signal output
rlabel metal3 s 59200 15784 60000 15904 6 s0_wbd_adr_o[14]
port 758 nsew signal output
rlabel metal3 s 59200 15512 60000 15632 6 s0_wbd_adr_o[15]
port 759 nsew signal output
rlabel metal3 s 59200 15240 60000 15360 6 s0_wbd_adr_o[16]
port 760 nsew signal output
rlabel metal3 s 59200 14968 60000 15088 6 s0_wbd_adr_o[17]
port 761 nsew signal output
rlabel metal3 s 59200 14696 60000 14816 6 s0_wbd_adr_o[18]
port 762 nsew signal output
rlabel metal3 s 59200 14424 60000 14544 6 s0_wbd_adr_o[19]
port 763 nsew signal output
rlabel metal3 s 59200 19320 60000 19440 6 s0_wbd_adr_o[1]
port 764 nsew signal output
rlabel metal3 s 59200 14152 60000 14272 6 s0_wbd_adr_o[20]
port 765 nsew signal output
rlabel metal3 s 59200 13880 60000 14000 6 s0_wbd_adr_o[21]
port 766 nsew signal output
rlabel metal3 s 59200 13608 60000 13728 6 s0_wbd_adr_o[22]
port 767 nsew signal output
rlabel metal3 s 59200 13336 60000 13456 6 s0_wbd_adr_o[23]
port 768 nsew signal output
rlabel metal3 s 59200 13064 60000 13184 6 s0_wbd_adr_o[24]
port 769 nsew signal output
rlabel metal3 s 59200 12792 60000 12912 6 s0_wbd_adr_o[25]
port 770 nsew signal output
rlabel metal3 s 59200 12520 60000 12640 6 s0_wbd_adr_o[26]
port 771 nsew signal output
rlabel metal3 s 59200 12248 60000 12368 6 s0_wbd_adr_o[27]
port 772 nsew signal output
rlabel metal3 s 59200 11976 60000 12096 6 s0_wbd_adr_o[28]
port 773 nsew signal output
rlabel metal3 s 59200 11704 60000 11824 6 s0_wbd_adr_o[29]
port 774 nsew signal output
rlabel metal3 s 59200 19048 60000 19168 6 s0_wbd_adr_o[2]
port 775 nsew signal output
rlabel metal3 s 59200 11432 60000 11552 6 s0_wbd_adr_o[30]
port 776 nsew signal output
rlabel metal3 s 59200 11160 60000 11280 6 s0_wbd_adr_o[31]
port 777 nsew signal output
rlabel metal3 s 59200 18776 60000 18896 6 s0_wbd_adr_o[3]
port 778 nsew signal output
rlabel metal3 s 59200 18504 60000 18624 6 s0_wbd_adr_o[4]
port 779 nsew signal output
rlabel metal3 s 59200 18232 60000 18352 6 s0_wbd_adr_o[5]
port 780 nsew signal output
rlabel metal3 s 59200 17960 60000 18080 6 s0_wbd_adr_o[6]
port 781 nsew signal output
rlabel metal3 s 59200 17688 60000 17808 6 s0_wbd_adr_o[7]
port 782 nsew signal output
rlabel metal3 s 59200 17416 60000 17536 6 s0_wbd_adr_o[8]
port 783 nsew signal output
rlabel metal3 s 59200 17144 60000 17264 6 s0_wbd_adr_o[9]
port 784 nsew signal output
rlabel metal3 s 59200 23400 60000 23520 6 s0_wbd_bl_o[0]
port 785 nsew signal output
rlabel metal3 s 59200 23128 60000 23248 6 s0_wbd_bl_o[1]
port 786 nsew signal output
rlabel metal3 s 59200 22856 60000 22976 6 s0_wbd_bl_o[2]
port 787 nsew signal output
rlabel metal3 s 59200 22584 60000 22704 6 s0_wbd_bl_o[3]
port 788 nsew signal output
rlabel metal3 s 59200 22312 60000 22432 6 s0_wbd_bl_o[4]
port 789 nsew signal output
rlabel metal3 s 59200 22040 60000 22160 6 s0_wbd_bl_o[5]
port 790 nsew signal output
rlabel metal3 s 59200 21768 60000 21888 6 s0_wbd_bl_o[6]
port 791 nsew signal output
rlabel metal3 s 59200 21496 60000 21616 6 s0_wbd_bl_o[7]
port 792 nsew signal output
rlabel metal3 s 59200 21224 60000 21344 6 s0_wbd_bl_o[8]
port 793 nsew signal output
rlabel metal3 s 59200 20952 60000 21072 6 s0_wbd_bl_o[9]
port 794 nsew signal output
rlabel metal3 s 59200 23672 60000 23792 6 s0_wbd_bry_o
port 795 nsew signal output
rlabel metal3 s 59200 41896 60000 42016 6 s0_wbd_cyc_o
port 796 nsew signal output
rlabel metal3 s 59200 41080 60000 41200 6 s0_wbd_dat_i[0]
port 797 nsew signal input
rlabel metal3 s 59200 38360 60000 38480 6 s0_wbd_dat_i[10]
port 798 nsew signal input
rlabel metal3 s 59200 38088 60000 38208 6 s0_wbd_dat_i[11]
port 799 nsew signal input
rlabel metal3 s 59200 37816 60000 37936 6 s0_wbd_dat_i[12]
port 800 nsew signal input
rlabel metal3 s 59200 37544 60000 37664 6 s0_wbd_dat_i[13]
port 801 nsew signal input
rlabel metal3 s 59200 37272 60000 37392 6 s0_wbd_dat_i[14]
port 802 nsew signal input
rlabel metal3 s 59200 37000 60000 37120 6 s0_wbd_dat_i[15]
port 803 nsew signal input
rlabel metal3 s 59200 36728 60000 36848 6 s0_wbd_dat_i[16]
port 804 nsew signal input
rlabel metal3 s 59200 36456 60000 36576 6 s0_wbd_dat_i[17]
port 805 nsew signal input
rlabel metal3 s 59200 36184 60000 36304 6 s0_wbd_dat_i[18]
port 806 nsew signal input
rlabel metal3 s 59200 35912 60000 36032 6 s0_wbd_dat_i[19]
port 807 nsew signal input
rlabel metal3 s 59200 40808 60000 40928 6 s0_wbd_dat_i[1]
port 808 nsew signal input
rlabel metal3 s 59200 35640 60000 35760 6 s0_wbd_dat_i[20]
port 809 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 s0_wbd_dat_i[21]
port 810 nsew signal input
rlabel metal3 s 59200 35096 60000 35216 6 s0_wbd_dat_i[22]
port 811 nsew signal input
rlabel metal3 s 59200 34824 60000 34944 6 s0_wbd_dat_i[23]
port 812 nsew signal input
rlabel metal3 s 59200 34552 60000 34672 6 s0_wbd_dat_i[24]
port 813 nsew signal input
rlabel metal3 s 59200 34280 60000 34400 6 s0_wbd_dat_i[25]
port 814 nsew signal input
rlabel metal3 s 59200 34008 60000 34128 6 s0_wbd_dat_i[26]
port 815 nsew signal input
rlabel metal3 s 59200 33736 60000 33856 6 s0_wbd_dat_i[27]
port 816 nsew signal input
rlabel metal3 s 59200 33464 60000 33584 6 s0_wbd_dat_i[28]
port 817 nsew signal input
rlabel metal3 s 59200 33192 60000 33312 6 s0_wbd_dat_i[29]
port 818 nsew signal input
rlabel metal3 s 59200 40536 60000 40656 6 s0_wbd_dat_i[2]
port 819 nsew signal input
rlabel metal3 s 59200 32920 60000 33040 6 s0_wbd_dat_i[30]
port 820 nsew signal input
rlabel metal3 s 59200 32648 60000 32768 6 s0_wbd_dat_i[31]
port 821 nsew signal input
rlabel metal3 s 59200 40264 60000 40384 6 s0_wbd_dat_i[3]
port 822 nsew signal input
rlabel metal3 s 59200 39992 60000 40112 6 s0_wbd_dat_i[4]
port 823 nsew signal input
rlabel metal3 s 59200 39720 60000 39840 6 s0_wbd_dat_i[5]
port 824 nsew signal input
rlabel metal3 s 59200 39448 60000 39568 6 s0_wbd_dat_i[6]
port 825 nsew signal input
rlabel metal3 s 59200 39176 60000 39296 6 s0_wbd_dat_i[7]
port 826 nsew signal input
rlabel metal3 s 59200 38904 60000 39024 6 s0_wbd_dat_i[8]
port 827 nsew signal input
rlabel metal3 s 59200 38632 60000 38752 6 s0_wbd_dat_i[9]
port 828 nsew signal input
rlabel metal3 s 59200 32376 60000 32496 6 s0_wbd_dat_o[0]
port 829 nsew signal output
rlabel metal3 s 59200 29656 60000 29776 6 s0_wbd_dat_o[10]
port 830 nsew signal output
rlabel metal3 s 59200 29384 60000 29504 6 s0_wbd_dat_o[11]
port 831 nsew signal output
rlabel metal3 s 59200 29112 60000 29232 6 s0_wbd_dat_o[12]
port 832 nsew signal output
rlabel metal3 s 59200 28840 60000 28960 6 s0_wbd_dat_o[13]
port 833 nsew signal output
rlabel metal3 s 59200 28568 60000 28688 6 s0_wbd_dat_o[14]
port 834 nsew signal output
rlabel metal3 s 59200 28296 60000 28416 6 s0_wbd_dat_o[15]
port 835 nsew signal output
rlabel metal3 s 59200 28024 60000 28144 6 s0_wbd_dat_o[16]
port 836 nsew signal output
rlabel metal3 s 59200 27752 60000 27872 6 s0_wbd_dat_o[17]
port 837 nsew signal output
rlabel metal3 s 59200 27480 60000 27600 6 s0_wbd_dat_o[18]
port 838 nsew signal output
rlabel metal3 s 59200 27208 60000 27328 6 s0_wbd_dat_o[19]
port 839 nsew signal output
rlabel metal3 s 59200 32104 60000 32224 6 s0_wbd_dat_o[1]
port 840 nsew signal output
rlabel metal3 s 59200 26936 60000 27056 6 s0_wbd_dat_o[20]
port 841 nsew signal output
rlabel metal3 s 59200 26664 60000 26784 6 s0_wbd_dat_o[21]
port 842 nsew signal output
rlabel metal3 s 59200 26392 60000 26512 6 s0_wbd_dat_o[22]
port 843 nsew signal output
rlabel metal3 s 59200 26120 60000 26240 6 s0_wbd_dat_o[23]
port 844 nsew signal output
rlabel metal3 s 59200 25848 60000 25968 6 s0_wbd_dat_o[24]
port 845 nsew signal output
rlabel metal3 s 59200 25576 60000 25696 6 s0_wbd_dat_o[25]
port 846 nsew signal output
rlabel metal3 s 59200 25304 60000 25424 6 s0_wbd_dat_o[26]
port 847 nsew signal output
rlabel metal3 s 59200 25032 60000 25152 6 s0_wbd_dat_o[27]
port 848 nsew signal output
rlabel metal3 s 59200 24760 60000 24880 6 s0_wbd_dat_o[28]
port 849 nsew signal output
rlabel metal3 s 59200 24488 60000 24608 6 s0_wbd_dat_o[29]
port 850 nsew signal output
rlabel metal3 s 59200 31832 60000 31952 6 s0_wbd_dat_o[2]
port 851 nsew signal output
rlabel metal3 s 59200 24216 60000 24336 6 s0_wbd_dat_o[30]
port 852 nsew signal output
rlabel metal3 s 59200 23944 60000 24064 6 s0_wbd_dat_o[31]
port 853 nsew signal output
rlabel metal3 s 59200 31560 60000 31680 6 s0_wbd_dat_o[3]
port 854 nsew signal output
rlabel metal3 s 59200 31288 60000 31408 6 s0_wbd_dat_o[4]
port 855 nsew signal output
rlabel metal3 s 59200 31016 60000 31136 6 s0_wbd_dat_o[5]
port 856 nsew signal output
rlabel metal3 s 59200 30744 60000 30864 6 s0_wbd_dat_o[6]
port 857 nsew signal output
rlabel metal3 s 59200 30472 60000 30592 6 s0_wbd_dat_o[7]
port 858 nsew signal output
rlabel metal3 s 59200 30200 60000 30320 6 s0_wbd_dat_o[8]
port 859 nsew signal output
rlabel metal3 s 59200 29928 60000 30048 6 s0_wbd_dat_o[9]
port 860 nsew signal output
rlabel metal3 s 59200 41624 60000 41744 6 s0_wbd_lack_i
port 861 nsew signal input
rlabel metal3 s 59200 20680 60000 20800 6 s0_wbd_sel_o[0]
port 862 nsew signal output
rlabel metal3 s 59200 20408 60000 20528 6 s0_wbd_sel_o[1]
port 863 nsew signal output
rlabel metal3 s 59200 20136 60000 20256 6 s0_wbd_sel_o[2]
port 864 nsew signal output
rlabel metal3 s 59200 19864 60000 19984 6 s0_wbd_sel_o[3]
port 865 nsew signal output
rlabel metal3 s 59200 10616 60000 10736 6 s0_wbd_stb_o
port 866 nsew signal output
rlabel metal3 s 59200 10888 60000 11008 6 s0_wbd_we_o
port 867 nsew signal output
rlabel metal3 s 59200 150016 60000 150136 6 s1_mclk
port 868 nsew signal output
rlabel metal3 s 59200 171776 60000 171896 6 s1_wbd_ack_i
port 869 nsew signal input
rlabel metal3 s 59200 153008 60000 153128 6 s1_wbd_adr_o[0]
port 870 nsew signal output
rlabel metal3 s 59200 152736 60000 152856 6 s1_wbd_adr_o[1]
port 871 nsew signal output
rlabel metal3 s 59200 152464 60000 152584 6 s1_wbd_adr_o[2]
port 872 nsew signal output
rlabel metal3 s 59200 152192 60000 152312 6 s1_wbd_adr_o[3]
port 873 nsew signal output
rlabel metal3 s 59200 151920 60000 152040 6 s1_wbd_adr_o[4]
port 874 nsew signal output
rlabel metal3 s 59200 151648 60000 151768 6 s1_wbd_adr_o[5]
port 875 nsew signal output
rlabel metal3 s 59200 151376 60000 151496 6 s1_wbd_adr_o[6]
port 876 nsew signal output
rlabel metal3 s 59200 151104 60000 151224 6 s1_wbd_adr_o[7]
port 877 nsew signal output
rlabel metal3 s 59200 150832 60000 150952 6 s1_wbd_adr_o[8]
port 878 nsew signal output
rlabel metal3 s 59200 172048 60000 172168 6 s1_wbd_cyc_o
port 879 nsew signal output
rlabel metal3 s 59200 171504 60000 171624 6 s1_wbd_dat_i[0]
port 880 nsew signal input
rlabel metal3 s 59200 168784 60000 168904 6 s1_wbd_dat_i[10]
port 881 nsew signal input
rlabel metal3 s 59200 168512 60000 168632 6 s1_wbd_dat_i[11]
port 882 nsew signal input
rlabel metal3 s 59200 168240 60000 168360 6 s1_wbd_dat_i[12]
port 883 nsew signal input
rlabel metal3 s 59200 167968 60000 168088 6 s1_wbd_dat_i[13]
port 884 nsew signal input
rlabel metal3 s 59200 167696 60000 167816 6 s1_wbd_dat_i[14]
port 885 nsew signal input
rlabel metal3 s 59200 167424 60000 167544 6 s1_wbd_dat_i[15]
port 886 nsew signal input
rlabel metal3 s 59200 167152 60000 167272 6 s1_wbd_dat_i[16]
port 887 nsew signal input
rlabel metal3 s 59200 166880 60000 167000 6 s1_wbd_dat_i[17]
port 888 nsew signal input
rlabel metal3 s 59200 166608 60000 166728 6 s1_wbd_dat_i[18]
port 889 nsew signal input
rlabel metal3 s 59200 166336 60000 166456 6 s1_wbd_dat_i[19]
port 890 nsew signal input
rlabel metal3 s 59200 171232 60000 171352 6 s1_wbd_dat_i[1]
port 891 nsew signal input
rlabel metal3 s 59200 166064 60000 166184 6 s1_wbd_dat_i[20]
port 892 nsew signal input
rlabel metal3 s 59200 165792 60000 165912 6 s1_wbd_dat_i[21]
port 893 nsew signal input
rlabel metal3 s 59200 165520 60000 165640 6 s1_wbd_dat_i[22]
port 894 nsew signal input
rlabel metal3 s 59200 165248 60000 165368 6 s1_wbd_dat_i[23]
port 895 nsew signal input
rlabel metal3 s 59200 164976 60000 165096 6 s1_wbd_dat_i[24]
port 896 nsew signal input
rlabel metal3 s 59200 164704 60000 164824 6 s1_wbd_dat_i[25]
port 897 nsew signal input
rlabel metal3 s 59200 164432 60000 164552 6 s1_wbd_dat_i[26]
port 898 nsew signal input
rlabel metal3 s 59200 164160 60000 164280 6 s1_wbd_dat_i[27]
port 899 nsew signal input
rlabel metal3 s 59200 163888 60000 164008 6 s1_wbd_dat_i[28]
port 900 nsew signal input
rlabel metal3 s 59200 163616 60000 163736 6 s1_wbd_dat_i[29]
port 901 nsew signal input
rlabel metal3 s 59200 170960 60000 171080 6 s1_wbd_dat_i[2]
port 902 nsew signal input
rlabel metal3 s 59200 163344 60000 163464 6 s1_wbd_dat_i[30]
port 903 nsew signal input
rlabel metal3 s 59200 163072 60000 163192 6 s1_wbd_dat_i[31]
port 904 nsew signal input
rlabel metal3 s 59200 170688 60000 170808 6 s1_wbd_dat_i[3]
port 905 nsew signal input
rlabel metal3 s 59200 170416 60000 170536 6 s1_wbd_dat_i[4]
port 906 nsew signal input
rlabel metal3 s 59200 170144 60000 170264 6 s1_wbd_dat_i[5]
port 907 nsew signal input
rlabel metal3 s 59200 169872 60000 169992 6 s1_wbd_dat_i[6]
port 908 nsew signal input
rlabel metal3 s 59200 169600 60000 169720 6 s1_wbd_dat_i[7]
port 909 nsew signal input
rlabel metal3 s 59200 169328 60000 169448 6 s1_wbd_dat_i[8]
port 910 nsew signal input
rlabel metal3 s 59200 169056 60000 169176 6 s1_wbd_dat_i[9]
port 911 nsew signal input
rlabel metal3 s 59200 162800 60000 162920 6 s1_wbd_dat_o[0]
port 912 nsew signal output
rlabel metal3 s 59200 160080 60000 160200 6 s1_wbd_dat_o[10]
port 913 nsew signal output
rlabel metal3 s 59200 159808 60000 159928 6 s1_wbd_dat_o[11]
port 914 nsew signal output
rlabel metal3 s 59200 159536 60000 159656 6 s1_wbd_dat_o[12]
port 915 nsew signal output
rlabel metal3 s 59200 159264 60000 159384 6 s1_wbd_dat_o[13]
port 916 nsew signal output
rlabel metal3 s 59200 158992 60000 159112 6 s1_wbd_dat_o[14]
port 917 nsew signal output
rlabel metal3 s 59200 158720 60000 158840 6 s1_wbd_dat_o[15]
port 918 nsew signal output
rlabel metal3 s 59200 158448 60000 158568 6 s1_wbd_dat_o[16]
port 919 nsew signal output
rlabel metal3 s 59200 158176 60000 158296 6 s1_wbd_dat_o[17]
port 920 nsew signal output
rlabel metal3 s 59200 157904 60000 158024 6 s1_wbd_dat_o[18]
port 921 nsew signal output
rlabel metal3 s 59200 157632 60000 157752 6 s1_wbd_dat_o[19]
port 922 nsew signal output
rlabel metal3 s 59200 162528 60000 162648 6 s1_wbd_dat_o[1]
port 923 nsew signal output
rlabel metal3 s 59200 157360 60000 157480 6 s1_wbd_dat_o[20]
port 924 nsew signal output
rlabel metal3 s 59200 157088 60000 157208 6 s1_wbd_dat_o[21]
port 925 nsew signal output
rlabel metal3 s 59200 156816 60000 156936 6 s1_wbd_dat_o[22]
port 926 nsew signal output
rlabel metal3 s 59200 156544 60000 156664 6 s1_wbd_dat_o[23]
port 927 nsew signal output
rlabel metal3 s 59200 156272 60000 156392 6 s1_wbd_dat_o[24]
port 928 nsew signal output
rlabel metal3 s 59200 156000 60000 156120 6 s1_wbd_dat_o[25]
port 929 nsew signal output
rlabel metal3 s 59200 155728 60000 155848 6 s1_wbd_dat_o[26]
port 930 nsew signal output
rlabel metal3 s 59200 155456 60000 155576 6 s1_wbd_dat_o[27]
port 931 nsew signal output
rlabel metal3 s 59200 155184 60000 155304 6 s1_wbd_dat_o[28]
port 932 nsew signal output
rlabel metal3 s 59200 154912 60000 155032 6 s1_wbd_dat_o[29]
port 933 nsew signal output
rlabel metal3 s 59200 162256 60000 162376 6 s1_wbd_dat_o[2]
port 934 nsew signal output
rlabel metal3 s 59200 154640 60000 154760 6 s1_wbd_dat_o[30]
port 935 nsew signal output
rlabel metal3 s 59200 154368 60000 154488 6 s1_wbd_dat_o[31]
port 936 nsew signal output
rlabel metal3 s 59200 161984 60000 162104 6 s1_wbd_dat_o[3]
port 937 nsew signal output
rlabel metal3 s 59200 161712 60000 161832 6 s1_wbd_dat_o[4]
port 938 nsew signal output
rlabel metal3 s 59200 161440 60000 161560 6 s1_wbd_dat_o[5]
port 939 nsew signal output
rlabel metal3 s 59200 161168 60000 161288 6 s1_wbd_dat_o[6]
port 940 nsew signal output
rlabel metal3 s 59200 160896 60000 161016 6 s1_wbd_dat_o[7]
port 941 nsew signal output
rlabel metal3 s 59200 160624 60000 160744 6 s1_wbd_dat_o[8]
port 942 nsew signal output
rlabel metal3 s 59200 160352 60000 160472 6 s1_wbd_dat_o[9]
port 943 nsew signal output
rlabel metal3 s 59200 154096 60000 154216 6 s1_wbd_sel_o[0]
port 944 nsew signal output
rlabel metal3 s 59200 153824 60000 153944 6 s1_wbd_sel_o[1]
port 945 nsew signal output
rlabel metal3 s 59200 153552 60000 153672 6 s1_wbd_sel_o[2]
port 946 nsew signal output
rlabel metal3 s 59200 153280 60000 153400 6 s1_wbd_sel_o[3]
port 947 nsew signal output
rlabel metal3 s 59200 150288 60000 150408 6 s1_wbd_stb_o
port 948 nsew signal output
rlabel metal3 s 59200 150560 60000 150680 6 s1_wbd_we_o
port 949 nsew signal output
rlabel metal3 s 59200 282072 60000 282192 6 s2_mclk
port 950 nsew signal output
rlabel metal3 s 59200 304376 60000 304496 6 s2_wbd_ack_i
port 951 nsew signal input
rlabel metal3 s 59200 285608 60000 285728 6 s2_wbd_adr_o[0]
port 952 nsew signal output
rlabel metal3 s 59200 282888 60000 283008 6 s2_wbd_adr_o[10]
port 953 nsew signal output
rlabel metal3 s 59200 285336 60000 285456 6 s2_wbd_adr_o[1]
port 954 nsew signal output
rlabel metal3 s 59200 285064 60000 285184 6 s2_wbd_adr_o[2]
port 955 nsew signal output
rlabel metal3 s 59200 284792 60000 284912 6 s2_wbd_adr_o[3]
port 956 nsew signal output
rlabel metal3 s 59200 284520 60000 284640 6 s2_wbd_adr_o[4]
port 957 nsew signal output
rlabel metal3 s 59200 284248 60000 284368 6 s2_wbd_adr_o[5]
port 958 nsew signal output
rlabel metal3 s 59200 283976 60000 284096 6 s2_wbd_adr_o[6]
port 959 nsew signal output
rlabel metal3 s 59200 283704 60000 283824 6 s2_wbd_adr_o[7]
port 960 nsew signal output
rlabel metal3 s 59200 283432 60000 283552 6 s2_wbd_adr_o[8]
port 961 nsew signal output
rlabel metal3 s 59200 283160 60000 283280 6 s2_wbd_adr_o[9]
port 962 nsew signal output
rlabel metal3 s 59200 304648 60000 304768 6 s2_wbd_cyc_o
port 963 nsew signal output
rlabel metal3 s 59200 304104 60000 304224 6 s2_wbd_dat_i[0]
port 964 nsew signal input
rlabel metal3 s 59200 301384 60000 301504 6 s2_wbd_dat_i[10]
port 965 nsew signal input
rlabel metal3 s 59200 301112 60000 301232 6 s2_wbd_dat_i[11]
port 966 nsew signal input
rlabel metal3 s 59200 300840 60000 300960 6 s2_wbd_dat_i[12]
port 967 nsew signal input
rlabel metal3 s 59200 300568 60000 300688 6 s2_wbd_dat_i[13]
port 968 nsew signal input
rlabel metal3 s 59200 300296 60000 300416 6 s2_wbd_dat_i[14]
port 969 nsew signal input
rlabel metal3 s 59200 300024 60000 300144 6 s2_wbd_dat_i[15]
port 970 nsew signal input
rlabel metal3 s 59200 299752 60000 299872 6 s2_wbd_dat_i[16]
port 971 nsew signal input
rlabel metal3 s 59200 299480 60000 299600 6 s2_wbd_dat_i[17]
port 972 nsew signal input
rlabel metal3 s 59200 299208 60000 299328 6 s2_wbd_dat_i[18]
port 973 nsew signal input
rlabel metal3 s 59200 298936 60000 299056 6 s2_wbd_dat_i[19]
port 974 nsew signal input
rlabel metal3 s 59200 303832 60000 303952 6 s2_wbd_dat_i[1]
port 975 nsew signal input
rlabel metal3 s 59200 298664 60000 298784 6 s2_wbd_dat_i[20]
port 976 nsew signal input
rlabel metal3 s 59200 298392 60000 298512 6 s2_wbd_dat_i[21]
port 977 nsew signal input
rlabel metal3 s 59200 298120 60000 298240 6 s2_wbd_dat_i[22]
port 978 nsew signal input
rlabel metal3 s 59200 297848 60000 297968 6 s2_wbd_dat_i[23]
port 979 nsew signal input
rlabel metal3 s 59200 297576 60000 297696 6 s2_wbd_dat_i[24]
port 980 nsew signal input
rlabel metal3 s 59200 297304 60000 297424 6 s2_wbd_dat_i[25]
port 981 nsew signal input
rlabel metal3 s 59200 297032 60000 297152 6 s2_wbd_dat_i[26]
port 982 nsew signal input
rlabel metal3 s 59200 296760 60000 296880 6 s2_wbd_dat_i[27]
port 983 nsew signal input
rlabel metal3 s 59200 296488 60000 296608 6 s2_wbd_dat_i[28]
port 984 nsew signal input
rlabel metal3 s 59200 296216 60000 296336 6 s2_wbd_dat_i[29]
port 985 nsew signal input
rlabel metal3 s 59200 303560 60000 303680 6 s2_wbd_dat_i[2]
port 986 nsew signal input
rlabel metal3 s 59200 295944 60000 296064 6 s2_wbd_dat_i[30]
port 987 nsew signal input
rlabel metal3 s 59200 295672 60000 295792 6 s2_wbd_dat_i[31]
port 988 nsew signal input
rlabel metal3 s 59200 303288 60000 303408 6 s2_wbd_dat_i[3]
port 989 nsew signal input
rlabel metal3 s 59200 303016 60000 303136 6 s2_wbd_dat_i[4]
port 990 nsew signal input
rlabel metal3 s 59200 302744 60000 302864 6 s2_wbd_dat_i[5]
port 991 nsew signal input
rlabel metal3 s 59200 302472 60000 302592 6 s2_wbd_dat_i[6]
port 992 nsew signal input
rlabel metal3 s 59200 302200 60000 302320 6 s2_wbd_dat_i[7]
port 993 nsew signal input
rlabel metal3 s 59200 301928 60000 302048 6 s2_wbd_dat_i[8]
port 994 nsew signal input
rlabel metal3 s 59200 301656 60000 301776 6 s2_wbd_dat_i[9]
port 995 nsew signal input
rlabel metal3 s 59200 295400 60000 295520 6 s2_wbd_dat_o[0]
port 996 nsew signal output
rlabel metal3 s 59200 292680 60000 292800 6 s2_wbd_dat_o[10]
port 997 nsew signal output
rlabel metal3 s 59200 292408 60000 292528 6 s2_wbd_dat_o[11]
port 998 nsew signal output
rlabel metal3 s 59200 292136 60000 292256 6 s2_wbd_dat_o[12]
port 999 nsew signal output
rlabel metal3 s 59200 291864 60000 291984 6 s2_wbd_dat_o[13]
port 1000 nsew signal output
rlabel metal3 s 59200 291592 60000 291712 6 s2_wbd_dat_o[14]
port 1001 nsew signal output
rlabel metal3 s 59200 291320 60000 291440 6 s2_wbd_dat_o[15]
port 1002 nsew signal output
rlabel metal3 s 59200 291048 60000 291168 6 s2_wbd_dat_o[16]
port 1003 nsew signal output
rlabel metal3 s 59200 290776 60000 290896 6 s2_wbd_dat_o[17]
port 1004 nsew signal output
rlabel metal3 s 59200 290504 60000 290624 6 s2_wbd_dat_o[18]
port 1005 nsew signal output
rlabel metal3 s 59200 290232 60000 290352 6 s2_wbd_dat_o[19]
port 1006 nsew signal output
rlabel metal3 s 59200 295128 60000 295248 6 s2_wbd_dat_o[1]
port 1007 nsew signal output
rlabel metal3 s 59200 289960 60000 290080 6 s2_wbd_dat_o[20]
port 1008 nsew signal output
rlabel metal3 s 59200 289688 60000 289808 6 s2_wbd_dat_o[21]
port 1009 nsew signal output
rlabel metal3 s 59200 289416 60000 289536 6 s2_wbd_dat_o[22]
port 1010 nsew signal output
rlabel metal3 s 59200 289144 60000 289264 6 s2_wbd_dat_o[23]
port 1011 nsew signal output
rlabel metal3 s 59200 288872 60000 288992 6 s2_wbd_dat_o[24]
port 1012 nsew signal output
rlabel metal3 s 59200 288600 60000 288720 6 s2_wbd_dat_o[25]
port 1013 nsew signal output
rlabel metal3 s 59200 288328 60000 288448 6 s2_wbd_dat_o[26]
port 1014 nsew signal output
rlabel metal3 s 59200 288056 60000 288176 6 s2_wbd_dat_o[27]
port 1015 nsew signal output
rlabel metal3 s 59200 287784 60000 287904 6 s2_wbd_dat_o[28]
port 1016 nsew signal output
rlabel metal3 s 59200 287512 60000 287632 6 s2_wbd_dat_o[29]
port 1017 nsew signal output
rlabel metal3 s 59200 294856 60000 294976 6 s2_wbd_dat_o[2]
port 1018 nsew signal output
rlabel metal3 s 59200 287240 60000 287360 6 s2_wbd_dat_o[30]
port 1019 nsew signal output
rlabel metal3 s 59200 286968 60000 287088 6 s2_wbd_dat_o[31]
port 1020 nsew signal output
rlabel metal3 s 59200 294584 60000 294704 6 s2_wbd_dat_o[3]
port 1021 nsew signal output
rlabel metal3 s 59200 294312 60000 294432 6 s2_wbd_dat_o[4]
port 1022 nsew signal output
rlabel metal3 s 59200 294040 60000 294160 6 s2_wbd_dat_o[5]
port 1023 nsew signal output
rlabel metal3 s 59200 293768 60000 293888 6 s2_wbd_dat_o[6]
port 1024 nsew signal output
rlabel metal3 s 59200 293496 60000 293616 6 s2_wbd_dat_o[7]
port 1025 nsew signal output
rlabel metal3 s 59200 293224 60000 293344 6 s2_wbd_dat_o[8]
port 1026 nsew signal output
rlabel metal3 s 59200 292952 60000 293072 6 s2_wbd_dat_o[9]
port 1027 nsew signal output
rlabel metal3 s 59200 286696 60000 286816 6 s2_wbd_sel_o[0]
port 1028 nsew signal output
rlabel metal3 s 59200 286424 60000 286544 6 s2_wbd_sel_o[1]
port 1029 nsew signal output
rlabel metal3 s 59200 286152 60000 286272 6 s2_wbd_sel_o[2]
port 1030 nsew signal output
rlabel metal3 s 59200 285880 60000 286000 6 s2_wbd_sel_o[3]
port 1031 nsew signal output
rlabel metal3 s 59200 282344 60000 282464 6 s2_wbd_stb_o
port 1032 nsew signal output
rlabel metal3 s 59200 282616 60000 282736 6 s2_wbd_we_o
port 1033 nsew signal output
rlabel metal4 s 3748 2128 4988 357456 6 vccd1
port 1034 nsew power bidirectional
rlabel metal4 s 23748 2128 24988 357456 6 vccd1
port 1034 nsew power bidirectional
rlabel metal4 s 43748 2128 44988 357456 6 vccd1
port 1034 nsew power bidirectional
rlabel metal4 s 13748 2128 14988 357456 6 vssd1
port 1035 nsew ground bidirectional
rlabel metal4 s 33748 2128 34988 357456 6 vssd1
port 1035 nsew ground bidirectional
rlabel metal4 s 53748 2128 54988 357456 6 vssd1
port 1035 nsew ground bidirectional
rlabel metal2 s 13266 0 13322 800 6 wbd_clk_int
port 1036 nsew signal input
rlabel metal2 s 13450 0 13506 800 6 wbd_clk_wi
port 1037 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60000 360000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 42759168
string GDS_FILE /home/lx/projects/caravel_env/caravel_usb_test/openlane/wb_interconnect/runs/wb_interconnect/results/signoff/wb_interconnect.magic.gds
string GDS_START 1263676
<< end >>

