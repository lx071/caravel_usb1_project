// This is the unpowered netlist.
module bus_rep_south (ch_in,
    ch_out);
 input [252:0] ch_in;
 output [252:0] ch_out;

 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net15;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net16;
 wire net160;
 wire net161;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[0].u_buf_A  (.DIODE(ch_in[0]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[100].u_buf_A  (.DIODE(ch_in[100]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[101].u_buf_A  (.DIODE(ch_in[101]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[102].u_buf_A  (.DIODE(net161));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[103].u_buf_A  (.DIODE(ch_in[103]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[104].u_buf_A  (.DIODE(ch_in[104]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[105].u_buf_A  (.DIODE(net160));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[106].u_buf_A  (.DIODE(ch_in[106]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[107].u_buf_A  (.DIODE(net159));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[108].u_buf_A  (.DIODE(ch_in[108]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[109].u_buf_A  (.DIODE(net158));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[10].u_buf_A  (.DIODE(ch_in[10]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[110].u_buf_A  (.DIODE(ch_in[110]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[111].u_buf_A  (.DIODE(net157));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[112].u_buf_A  (.DIODE(ch_in[112]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[113].u_buf_A  (.DIODE(net156));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[114].u_buf_A  (.DIODE(ch_in[114]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[115].u_buf_A  (.DIODE(net155));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[116].u_buf_A  (.DIODE(ch_in[116]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[117].u_buf_A  (.DIODE(net154));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[118].u_buf_A  (.DIODE(ch_in[118]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[119].u_buf_A  (.DIODE(net153));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[11].u_buf_A  (.DIODE(ch_in[11]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[120].u_buf_A  (.DIODE(ch_in[120]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[121].u_buf_A  (.DIODE(net152));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[122].u_buf_A  (.DIODE(ch_in[122]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[123].u_buf_A  (.DIODE(net151));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[124].u_buf_A  (.DIODE(ch_in[124]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[125].u_buf_A  (.DIODE(net150));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[126].u_buf_A  (.DIODE(ch_in[126]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[127].u_buf_A  (.DIODE(net149));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[128].u_buf_A  (.DIODE(ch_in[128]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[129].u_buf_A  (.DIODE(net148));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[12].u_buf_A  (.DIODE(net147));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[130].u_buf_A  (.DIODE(ch_in[130]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[131].u_buf_A  (.DIODE(net146));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[132].u_buf_A  (.DIODE(ch_in[132]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[133].u_buf_A  (.DIODE(net145));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[134].u_buf_A  (.DIODE(ch_in[134]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[135].u_buf_A  (.DIODE(net144));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[136].u_buf_A  (.DIODE(ch_in[136]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[137].u_buf_A  (.DIODE(net143));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[138].u_buf_A  (.DIODE(ch_in[138]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[139].u_buf_A  (.DIODE(net142));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[13].u_buf_A  (.DIODE(ch_in[13]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[140].u_buf_A  (.DIODE(ch_in[140]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[141].u_buf_A  (.DIODE(net141));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[142].u_buf_A  (.DIODE(net140));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[143].u_buf_A  (.DIODE(net139));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[144].u_buf_A  (.DIODE(net138));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[145].u_buf_A  (.DIODE(net137));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[146].u_buf_A  (.DIODE(net136));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[147].u_buf_A  (.DIODE(net135));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[148].u_buf_A  (.DIODE(net134));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[149].u_buf_A  (.DIODE(net133));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[14].u_buf_A  (.DIODE(ch_in[14]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[150].u_buf_A  (.DIODE(net132));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[151].u_buf_A  (.DIODE(net131));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[152].u_buf_A  (.DIODE(net130));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[153].u_buf_A  (.DIODE(net129));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[154].u_buf_A  (.DIODE(net128));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[155].u_buf_A  (.DIODE(net127));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[156].u_buf_A  (.DIODE(net126));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[157].u_buf_A  (.DIODE(net125));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[158].u_buf_A  (.DIODE(net124));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[159].u_buf_A  (.DIODE(net123));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[15].u_buf_A  (.DIODE(ch_in[15]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[160].u_buf_A  (.DIODE(net122));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[161].u_buf_A  (.DIODE(ch_in[161]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[162].u_buf_A  (.DIODE(ch_in[162]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[163].u_buf_A  (.DIODE(ch_in[163]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[164].u_buf_A  (.DIODE(ch_in[164]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[165].u_buf_A  (.DIODE(ch_in[165]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[166].u_buf_A  (.DIODE(ch_in[166]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[167].u_buf_A  (.DIODE(ch_in[167]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[168].u_buf_A  (.DIODE(ch_in[168]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[169].u_buf_A  (.DIODE(ch_in[169]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[16].u_buf_A  (.DIODE(net121));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[170].u_buf_A  (.DIODE(ch_in[170]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[171].u_buf_A  (.DIODE(ch_in[171]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[172].u_buf_A  (.DIODE(ch_in[172]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[173].u_buf_A  (.DIODE(ch_in[173]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[174].u_buf_A  (.DIODE(ch_in[174]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[175].u_buf_A  (.DIODE(ch_in[175]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[176].u_buf_A  (.DIODE(ch_in[176]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[177].u_buf_A  (.DIODE(ch_in[177]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[178].u_buf_A  (.DIODE(ch_in[178]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[179].u_buf_A  (.DIODE(ch_in[179]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[17].u_buf_A  (.DIODE(ch_in[17]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[180].u_buf_A  (.DIODE(ch_in[180]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[181].u_buf_A  (.DIODE(ch_in[181]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[182].u_buf_A  (.DIODE(ch_in[182]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[183].u_buf_A  (.DIODE(ch_in[183]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[184].u_buf_A  (.DIODE(ch_in[184]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[185].u_buf_A  (.DIODE(ch_in[185]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[186].u_buf_A  (.DIODE(ch_in[186]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[187].u_buf_A  (.DIODE(ch_in[187]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[188].u_buf_A  (.DIODE(ch_in[188]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[189].u_buf_A  (.DIODE(ch_in[189]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[18].u_buf_A  (.DIODE(ch_in[18]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[190].u_buf_A  (.DIODE(ch_in[190]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[191].u_buf_A  (.DIODE(ch_in[191]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[192].u_buf_A  (.DIODE(ch_in[192]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[193].u_buf_A  (.DIODE(ch_in[193]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[194].u_buf_A  (.DIODE(ch_in[194]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[195].u_buf_A  (.DIODE(ch_in[195]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[196].u_buf_A  (.DIODE(ch_in[196]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[197].u_buf_A  (.DIODE(ch_in[197]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[198].u_buf_A  (.DIODE(ch_in[198]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[199].u_buf_A  (.DIODE(ch_in[199]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[19].u_buf_A  (.DIODE(ch_in[19]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[1].u_buf_A  (.DIODE(ch_in[1]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[200].u_buf_A  (.DIODE(ch_in[200]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[201].u_buf_A  (.DIODE(ch_in[201]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[202].u_buf_A  (.DIODE(ch_in[202]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[203].u_buf_A  (.DIODE(ch_in[203]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[204].u_buf_A  (.DIODE(ch_in[204]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[205].u_buf_A  (.DIODE(ch_in[205]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[206].u_buf_A  (.DIODE(ch_in[206]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[207].u_buf_A  (.DIODE(ch_in[207]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[208].u_buf_A  (.DIODE(ch_in[208]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[209].u_buf_A  (.DIODE(ch_in[209]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[20].u_buf_A  (.DIODE(net120));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[210].u_buf_A  (.DIODE(ch_in[210]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[211].u_buf_A  (.DIODE(ch_in[211]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[212].u_buf_A  (.DIODE(ch_in[212]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[213].u_buf_A  (.DIODE(ch_in[213]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[214].u_buf_A  (.DIODE(ch_in[214]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[215].u_buf_A  (.DIODE(ch_in[215]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[216].u_buf_A  (.DIODE(ch_in[216]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[217].u_buf_A  (.DIODE(ch_in[217]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[218].u_buf_A  (.DIODE(ch_in[218]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[219].u_buf_A  (.DIODE(ch_in[219]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[21].u_buf_A  (.DIODE(ch_in[21]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[220].u_buf_A  (.DIODE(ch_in[220]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[221].u_buf_A  (.DIODE(ch_in[221]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[222].u_buf_A  (.DIODE(ch_in[222]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[223].u_buf_A  (.DIODE(ch_in[223]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[224].u_buf_A  (.DIODE(ch_in[224]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[225].u_buf_A  (.DIODE(ch_in[225]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[226].u_buf_A  (.DIODE(ch_in[226]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[227].u_buf_A  (.DIODE(ch_in[227]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[228].u_buf_A  (.DIODE(ch_in[228]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[229].u_buf_A  (.DIODE(ch_in[229]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[22].u_buf_A  (.DIODE(ch_in[22]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[230].u_buf_A  (.DIODE(ch_in[230]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[231].u_buf_A  (.DIODE(ch_in[231]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[232].u_buf_A  (.DIODE(ch_in[232]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[233].u_buf_A  (.DIODE(ch_in[233]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[234].u_buf_A  (.DIODE(ch_in[234]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[235].u_buf_A  (.DIODE(ch_in[235]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[236].u_buf_A  (.DIODE(ch_in[236]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[237].u_buf_A  (.DIODE(ch_in[237]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[238].u_buf_A  (.DIODE(ch_in[238]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[239].u_buf_A  (.DIODE(ch_in[239]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[23].u_buf_A  (.DIODE(ch_in[23]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[240].u_buf_A  (.DIODE(ch_in[240]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[241].u_buf_A  (.DIODE(ch_in[241]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[242].u_buf_A  (.DIODE(ch_in[242]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[243].u_buf_A  (.DIODE(ch_in[243]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[244].u_buf_A  (.DIODE(ch_in[244]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[245].u_buf_A  (.DIODE(ch_in[245]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[246].u_buf_A  (.DIODE(ch_in[246]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[247].u_buf_A  (.DIODE(ch_in[247]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[248].u_buf_A  (.DIODE(ch_in[248]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[249].u_buf_A  (.DIODE(ch_in[249]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[24].u_buf_A  (.DIODE(net119));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[250].u_buf_A  (.DIODE(ch_in[250]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[251].u_buf_A  (.DIODE(ch_in[251]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[252].u_buf_A  (.DIODE(ch_in[252]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[25].u_buf_A  (.DIODE(ch_in[25]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[26].u_buf_A  (.DIODE(ch_in[26]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[27].u_buf_A  (.DIODE(net118));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[28].u_buf_A  (.DIODE(ch_in[28]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[29].u_buf_A  (.DIODE(ch_in[29]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[2].u_buf_A  (.DIODE(net117));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[30].u_buf_A  (.DIODE(net116));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[31].u_buf_A  (.DIODE(ch_in[31]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[32].u_buf_A  (.DIODE(ch_in[32]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[33].u_buf_A  (.DIODE(net115));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[34].u_buf_A  (.DIODE(ch_in[34]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[35].u_buf_A  (.DIODE(ch_in[35]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[36].u_buf_A  (.DIODE(net114));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[37].u_buf_A  (.DIODE(ch_in[37]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[38].u_buf_A  (.DIODE(ch_in[38]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[39].u_buf_A  (.DIODE(net113));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[3].u_buf_A  (.DIODE(ch_in[3]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[40].u_buf_A  (.DIODE(ch_in[40]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[41].u_buf_A  (.DIODE(ch_in[41]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[42].u_buf_A  (.DIODE(net112));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[43].u_buf_A  (.DIODE(ch_in[43]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[44].u_buf_A  (.DIODE(ch_in[44]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[45].u_buf_A  (.DIODE(net111));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[46].u_buf_A  (.DIODE(ch_in[46]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[47].u_buf_A  (.DIODE(ch_in[47]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[48].u_buf_A  (.DIODE(net110));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[49].u_buf_A  (.DIODE(ch_in[49]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[4].u_buf_A  (.DIODE(ch_in[4]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[50].u_buf_A  (.DIODE(ch_in[50]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[51].u_buf_A  (.DIODE(net109));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[52].u_buf_A  (.DIODE(ch_in[52]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[53].u_buf_A  (.DIODE(ch_in[53]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[54].u_buf_A  (.DIODE(net108));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[55].u_buf_A  (.DIODE(ch_in[55]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[56].u_buf_A  (.DIODE(ch_in[56]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[57].u_buf_A  (.DIODE(net107));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[58].u_buf_A  (.DIODE(ch_in[58]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[59].u_buf_A  (.DIODE(ch_in[59]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[5].u_buf_A  (.DIODE(ch_in[5]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[60].u_buf_A  (.DIODE(net106));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[61].u_buf_A  (.DIODE(ch_in[61]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[62].u_buf_A  (.DIODE(ch_in[62]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[63].u_buf_A  (.DIODE(net105));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[64].u_buf_A  (.DIODE(ch_in[64]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[65].u_buf_A  (.DIODE(ch_in[65]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[66].u_buf_A  (.DIODE(net104));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[67].u_buf_A  (.DIODE(ch_in[67]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[68].u_buf_A  (.DIODE(ch_in[68]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[69].u_buf_A  (.DIODE(net103));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[6].u_buf_A  (.DIODE(ch_in[6]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[70].u_buf_A  (.DIODE(ch_in[70]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[71].u_buf_A  (.DIODE(ch_in[71]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[72].u_buf_A  (.DIODE(net102));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[73].u_buf_A  (.DIODE(ch_in[73]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[74].u_buf_A  (.DIODE(ch_in[74]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[75].u_buf_A  (.DIODE(net101));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[76].u_buf_A  (.DIODE(ch_in[76]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[77].u_buf_A  (.DIODE(ch_in[77]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[78].u_buf_A  (.DIODE(net100));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[79].u_buf_A  (.DIODE(ch_in[79]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[7].u_buf_A  (.DIODE(ch_in[7]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[80].u_buf_A  (.DIODE(ch_in[80]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[81].u_buf_A  (.DIODE(net99));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[82].u_buf_A  (.DIODE(ch_in[82]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[83].u_buf_A  (.DIODE(ch_in[83]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[84].u_buf_A  (.DIODE(net98));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[85].u_buf_A  (.DIODE(ch_in[85]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[86].u_buf_A  (.DIODE(ch_in[86]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[87].u_buf_A  (.DIODE(net97));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[88].u_buf_A  (.DIODE(ch_in[88]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[89].u_buf_A  (.DIODE(ch_in[89]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[8].u_buf_A  (.DIODE(net96));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[90].u_buf_A  (.DIODE(net95));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[91].u_buf_A  (.DIODE(ch_in[91]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[92].u_buf_A  (.DIODE(ch_in[92]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[93].u_buf_A  (.DIODE(net94));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[94].u_buf_A  (.DIODE(ch_in[94]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[95].u_buf_A  (.DIODE(ch_in[95]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[96].u_buf_A  (.DIODE(net93));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[97].u_buf_A  (.DIODE(ch_in[97]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[98].u_buf_A  (.DIODE(ch_in[98]));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[99].u_buf_A  (.DIODE(net92));
 sky130_fd_sc_hd__diode_2 \ANTENNA_u_rp[9].u_buf_A  (.DIODE(ch_in[9]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire100_A (.DIODE(ch_in[78]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire101_A (.DIODE(ch_in[75]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire102_A (.DIODE(ch_in[72]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire103_A (.DIODE(ch_in[69]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire104_A (.DIODE(ch_in[66]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire105_A (.DIODE(ch_in[63]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire106_A (.DIODE(ch_in[60]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire107_A (.DIODE(ch_in[57]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire108_A (.DIODE(ch_in[54]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire109_A (.DIODE(ch_in[51]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire10_A (.DIODE(net10));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire110_A (.DIODE(ch_in[48]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire111_A (.DIODE(ch_in[45]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire112_A (.DIODE(ch_in[42]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire113_A (.DIODE(ch_in[39]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire114_A (.DIODE(ch_in[36]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire115_A (.DIODE(ch_in[33]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire116_A (.DIODE(ch_in[30]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire117_A (.DIODE(ch_in[2]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire118_A (.DIODE(ch_in[27]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire119_A (.DIODE(ch_in[24]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire11_A (.DIODE(net11));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire120_A (.DIODE(ch_in[20]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire121_A (.DIODE(ch_in[16]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire122_A (.DIODE(ch_in[160]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire123_A (.DIODE(ch_in[159]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire124_A (.DIODE(ch_in[158]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire125_A (.DIODE(ch_in[157]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire126_A (.DIODE(ch_in[156]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire127_A (.DIODE(ch_in[155]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire128_A (.DIODE(ch_in[154]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire129_A (.DIODE(ch_in[153]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire12_A (.DIODE(net12));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire130_A (.DIODE(ch_in[152]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire131_A (.DIODE(ch_in[151]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire132_A (.DIODE(ch_in[150]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire133_A (.DIODE(ch_in[149]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire134_A (.DIODE(ch_in[148]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire135_A (.DIODE(ch_in[147]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire136_A (.DIODE(ch_in[146]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire137_A (.DIODE(ch_in[145]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire138_A (.DIODE(ch_in[144]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire139_A (.DIODE(ch_in[143]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire13_A (.DIODE(net13));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire140_A (.DIODE(ch_in[142]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire141_A (.DIODE(ch_in[141]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire142_A (.DIODE(ch_in[139]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire143_A (.DIODE(ch_in[137]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire144_A (.DIODE(ch_in[135]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire145_A (.DIODE(ch_in[133]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire146_A (.DIODE(ch_in[131]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire147_A (.DIODE(ch_in[12]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire148_A (.DIODE(ch_in[129]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire149_A (.DIODE(ch_in[127]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire14_A (.DIODE(net14));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire150_A (.DIODE(ch_in[125]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire151_A (.DIODE(ch_in[123]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire152_A (.DIODE(ch_in[121]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire153_A (.DIODE(ch_in[119]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire154_A (.DIODE(ch_in[117]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire155_A (.DIODE(ch_in[115]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire156_A (.DIODE(ch_in[113]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire157_A (.DIODE(ch_in[111]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire158_A (.DIODE(ch_in[109]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire159_A (.DIODE(ch_in[107]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire15_A (.DIODE(net15));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire160_A (.DIODE(ch_in[105]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire161_A (.DIODE(ch_in[102]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire16_A (.DIODE(net16));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire17_A (.DIODE(net17));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire18_A (.DIODE(net18));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire19_A (.DIODE(net19));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire1_A (.DIODE(net1));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire20_A (.DIODE(net20));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire21_A (.DIODE(net21));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire22_A (.DIODE(net22));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire23_A (.DIODE(net23));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire24_A (.DIODE(net24));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire25_A (.DIODE(net25));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire26_A (.DIODE(net26));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire27_A (.DIODE(net27));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire28_A (.DIODE(net28));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire29_A (.DIODE(net29));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire2_A (.DIODE(net2));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire30_A (.DIODE(net30));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire31_A (.DIODE(net31));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire32_A (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire33_A (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire34_A (.DIODE(net34));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire35_A (.DIODE(net35));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire36_A (.DIODE(net36));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire37_A (.DIODE(net37));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire38_A (.DIODE(net38));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire39_A (.DIODE(net39));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire3_A (.DIODE(net3));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire40_A (.DIODE(net40));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire41_A (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire42_A (.DIODE(net42));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire43_A (.DIODE(net43));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire44_A (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire45_A (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire46_A (.DIODE(net46));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire47_A (.DIODE(net47));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire48_A (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire49_A (.DIODE(net49));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire4_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire50_A (.DIODE(net50));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire51_A (.DIODE(net51));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire52_A (.DIODE(net52));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire53_A (.DIODE(net53));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire54_A (.DIODE(net54));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire55_A (.DIODE(net55));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire56_A (.DIODE(net56));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire57_A (.DIODE(net57));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire58_A (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire59_A (.DIODE(net59));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire5_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire60_A (.DIODE(net60));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire61_A (.DIODE(net61));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire62_A (.DIODE(net62));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire63_A (.DIODE(net63));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire64_A (.DIODE(net64));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire65_A (.DIODE(net65));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire66_A (.DIODE(net66));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire67_A (.DIODE(net67));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire68_A (.DIODE(net68));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire69_A (.DIODE(net69));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire6_A (.DIODE(net6));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire70_A (.DIODE(net70));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire71_A (.DIODE(net71));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire72_A (.DIODE(net72));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire73_A (.DIODE(net73));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire74_A (.DIODE(net74));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire75_A (.DIODE(net75));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire76_A (.DIODE(net76));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire77_A (.DIODE(net77));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire78_A (.DIODE(net78));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire79_A (.DIODE(net79));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire7_A (.DIODE(net7));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire80_A (.DIODE(net80));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire81_A (.DIODE(net81));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire82_A (.DIODE(net82));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire83_A (.DIODE(net83));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire84_A (.DIODE(net84));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire85_A (.DIODE(net85));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire86_A (.DIODE(net86));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire89_A (.DIODE(net89));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire8_A (.DIODE(net8));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire90_A (.DIODE(net90));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire91_A (.DIODE(net91));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire92_A (.DIODE(ch_in[99]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire93_A (.DIODE(ch_in[96]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire94_A (.DIODE(ch_in[93]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire95_A (.DIODE(ch_in[90]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire96_A (.DIODE(ch_in[8]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire97_A (.DIODE(ch_in[87]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire98_A (.DIODE(ch_in[84]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire99_A (.DIODE(ch_in[81]));
 sky130_fd_sc_hd__diode_2 ANTENNA_wire9_A (.DIODE(net9));
 sky130_fd_sc_hd__decap_4 FILLER_0_1003 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1007 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1019 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1033 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1047 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1059 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1063 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1103 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1143 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1159 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1227 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1261 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1271 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1285 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1299 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1314 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1327 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1343 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1361 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1399 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1463 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1495 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1511 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1579 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1623 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_163 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1635 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1679 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1691 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1697 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1705 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1719 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1731 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1735 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1737 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1775 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1787 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1791 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1793 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1803 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1831 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1843 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1847 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1849 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1859 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1865 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1887 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1899 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1903 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1905 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_191 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1915 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1921 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1933 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1943 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1955 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1959 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1961 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1971 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1977 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1999 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2011 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2015 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2017 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2027 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2033 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2041 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2055 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2067 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2071 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2073 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2083 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2123 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2127 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2145 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2179 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2183 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_219 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2201 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2241 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2265 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2279 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2295 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2351 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2369 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2407 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_247 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2509 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2573 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2587 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2605 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2621 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2649 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2661 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2689 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2733 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2741 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2783 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2789 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2797 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2801 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2811 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2817 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2825 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2829 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2839 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2845 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2853 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2867 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2873 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2881 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2885 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2901 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2909 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2913 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2923 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2929 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2937 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2941 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2951 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2957 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2965 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2969 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2979 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2985 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2993 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2997 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3007 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3013 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3021 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3025 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3035 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3041 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3049 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3053 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3063 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3069 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3077 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3081 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3091 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3097 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3105 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3137 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3147 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3217 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3245 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3259 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3273 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3329 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_335 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3389 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3413 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3441 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3473 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3497 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3529 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3539 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3557 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3581 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3585 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3613 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3637 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3641 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3735 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3763 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3777 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3791 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3805 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3819 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3833 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3847 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3861 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3875 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3889 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3893 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3903 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3909 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3917 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3921 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3931 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3945 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3949 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3959 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3965 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3973 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3977 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3987 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3993 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4001 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4005 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4015 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4033 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4043 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4057 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4061 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4071 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4085 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4089 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4099 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4117 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4145 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4173 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4183 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_419 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4201 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4211 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4217 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4239 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4245 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4267 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4285 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4295 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4313 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4323 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4329 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_437 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4379 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4393 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4397 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4413 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4435 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4453 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4463 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4491 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4497 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4519 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4547 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4565 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4575 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4603 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4617 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4621 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4631 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4637 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4649 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4659 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4665 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4677 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4693 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4715 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4721 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4733 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_474 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4743 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4749 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4761 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4777 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4785 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4789 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4799 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4805 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4813 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4817 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4827 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4833 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4841 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4845 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4855 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4861 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4873 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4883 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4889 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4897 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4901 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4911 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4917 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4925 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4929 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4939 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4945 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4953 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4957 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4967 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4973 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4981 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4985 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4995 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5001 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5009 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5013 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5023 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5029 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5037 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5041 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5051 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5057 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5065 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5069 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5079 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5085 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5093 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5163 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5191 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_521 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5275 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5287 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5291 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5303 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5315 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5331 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5347 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5387 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5399 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5403 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5431 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5443 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5455 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5471 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5487 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5499 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5511 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5527 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5543 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5555 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5571 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_613 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_627 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_642 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_671 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_767 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_773 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_781 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_785 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_795 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_807 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_810 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_813 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_823 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_835 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_839 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_841 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_851 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_857 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_865 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_879 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_891 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_895 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_925 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_935 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_941 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_963 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_975 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_978 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_991 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1007 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1012 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1020 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1025 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1033 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1041 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1051 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1063 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1075 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1083 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1088 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_121 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1217 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1221 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1237 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1249 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1285 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1297 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1314 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1321 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1345 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1369 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1413 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1424 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1433 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1457 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_1479 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1483 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1597 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1619 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1631 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_1643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2717 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2721 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_2965 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_2977 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2994 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3001 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3013 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3025 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3037 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3050 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3057 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3069 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3093 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3106 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3113 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3125 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3137 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3161 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3169 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3181 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3193 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_3215 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3219 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3225 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3237 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_979 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_986 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1534 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1540 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1552 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1585 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1597 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1679 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_1681 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1689 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1699 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1761 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1782 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_1788 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3249 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3270 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3276 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3288 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3300 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3305 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_3313 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3343 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3355 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3359 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3379 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3415 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3417 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_3434 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3440 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3452 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_3464 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1621 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_1633 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1650 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1709 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1721 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1734 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1740 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1752 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1789 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1801 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1807 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1817 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1825 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1837 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1849 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1864 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_1870 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1877 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_189 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1899 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_1929 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1933 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_1946 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1952 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1964 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1976 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2001 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2013 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2019 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2029 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_2035 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2585 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_2599 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3457 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3469 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_3477 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3488 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3494 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3513 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3525 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3533 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3543 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3587 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3597 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3603 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_3651 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_3657 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4027 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4039 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_4051 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_993 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1161 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1189 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1217 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1273 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1301 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1329 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1369 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1385 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1413 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1441 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1469 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1553 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1581 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1609 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1665 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1693 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1721 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1749 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1777 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1833 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1861 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1889 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1917 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1929 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1945 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_1982 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2005 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2029 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2041 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2045 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2053 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2064 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2070 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2097 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2101 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2112 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2118 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2126 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2129 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2146 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2152 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2169 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2181 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2185 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2196 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2202 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2210 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2213 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2225 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2253 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2265 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2269 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2277 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2283 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2295 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2297 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2307 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2313 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2337 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2349 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2353 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2367 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2379 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2381 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2395 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2409 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2421 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2427 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2434 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2441 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2453 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2461 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2465 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2479 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2493 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2509 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2516 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_2537 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2545 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2549 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2563 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2577 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2589 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2617 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2629 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_2633 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2647 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2673 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2689 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2701 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2729 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2757 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2785 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2813 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2841 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2869 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2953 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2981 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3009 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3037 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3049 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3065 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3093 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3121 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3149 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3177 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3233 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3261 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3289 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3317 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3329 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3345 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3373 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3401 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3429 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3457 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3513 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3541 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3569 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3597 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3609 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3625 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3653 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3665 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3669 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3680 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3686 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3694 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3697 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3708 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3714 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3722 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3725 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3736 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3742 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3750 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3753 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3767 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3779 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3781 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3789 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3795 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3807 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3809 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3823 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3835 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3837 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3845 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3851 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3863 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3865 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3873 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3879 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3883 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_389 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3890 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3897 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3909 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3918 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3937 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3945 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3953 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_3971 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_3975 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_3977 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_3981 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_3989 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_3998 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4005 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4009 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_4017 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4051 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4057 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4061 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4069 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4078 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4084 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4089 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4104 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4110 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4117 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4131 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4143 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_4145 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_4157 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_4163 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4185 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4213 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4241 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4269 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4297 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4353 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4381 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4409 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4437 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4449 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4465 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4493 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4521 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4549 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4577 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4633 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4661 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4689 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4717 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4729 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4745 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4773 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4801 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4829 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4857 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4913 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4941 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4969 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_4997 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5009 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5025 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5053 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5081 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5097 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5109 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5137 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5193 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5221 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5249 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5277 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5289 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5293 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5305 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5333 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5361 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5389 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5417 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5473 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5489 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5501 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5529 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5557 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5569 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5585 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5613 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5641 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5669 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_993 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1009 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1021 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1043 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1055 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1063 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1071 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1083 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1095 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1099 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1111 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1119 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1127 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1139 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1151 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1155 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1167 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1189 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1211 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1223 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1231 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1239 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1251 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1267 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1279 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1287 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1307 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_1319 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1323 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1335 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1357 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1369 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1391 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1469 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1489 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1525 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1545 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1557 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1569 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1581 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1601 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1613 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1637 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1649 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1669 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1693 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1713 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1725 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1749 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1769 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1781 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1825 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1837 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1861 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1881 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1893 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_19 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1917 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1929 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1937 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_1949 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1973 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_1993 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2005 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_201 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2029 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2049 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2061 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2085 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2105 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2117 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2129 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2141 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2163 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2175 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2197 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2209 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2219 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2231 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2253 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2275 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2287 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2309 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2331 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2343 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2387 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2399 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2421 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2443 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_2455 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2489 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2569 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2689 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2769 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2781 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_2993 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3049 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3129 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_313 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3249 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3297 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3329 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3341 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3609 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3689 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3809 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3889 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3901 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3921 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_3969 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4201 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4381 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4481 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4493 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4785 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4941 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5097 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5263 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5271 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5283 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5295 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5299 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5311 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5319 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5327 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5339 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5351 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5355 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5367 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5375 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5383 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_539 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5395 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5407 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5411 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5423 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5431 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5439 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5451 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5463 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5467 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5479 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5487 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5489 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5495 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5507 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_551 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5519 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5523 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5535 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5543 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5551 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5563 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_5575 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5579 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5591 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5601 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5693 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_607 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_635 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_727 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_735 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_747 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_759 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_763 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_775 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_783 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_791 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_803 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_815 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_819 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_831 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_841 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_853 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_875 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_887 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_89 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_895 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_903 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_915 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_927 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_931 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_943 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_951 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_959 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_971 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_983 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_987 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_999 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1003 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1019 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1031 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1035 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1037 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1047 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1053 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1067 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1075 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1087 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1091 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1103 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1115 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1131 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1137 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1145 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1159 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1171 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1179 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1187 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1199 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1203 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1205 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1215 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1235 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1243 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1255 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1259 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1271 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1283 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1305 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1327 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1339 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1347 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1355 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1367 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1371 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1373 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1383 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1401 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1407 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1411 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1417 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1425 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1429 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1435 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1439 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1445 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1457 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_1467 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_1473 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1521 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1595 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1601 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1625 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1637 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1689 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1889 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1901 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1969 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2081 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2181 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_219 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2205 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2249 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2293 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2449 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2461 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2529 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2641 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2741 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_275 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2765 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2809 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2897 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_2997 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3009 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3021 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3089 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_319 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3201 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3301 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3325 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3369 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_347 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3569 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3581 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3649 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3749 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3761 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3805 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3885 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3929 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_393 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4097 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4129 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4141 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4209 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_431 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4321 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4445 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4589 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4645 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4689 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4725 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4745 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4769 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_487 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4881 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4981 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5005 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5069 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5093 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5261 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5329 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5429 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5441 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5565 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5629 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5697 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_5721 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_599 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_667 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_699 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_711 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_717 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_731 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_755 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_779 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_795 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_801 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_809 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_823 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_835 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_843 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_851 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_863 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_867 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_869 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_879 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_885 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_899 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_907 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_919 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_923 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_935 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_947 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_963 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_969 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_977 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_991 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1469 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1487 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1499 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1511 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1524 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1536 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1546 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1556 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1566 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1569 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1577 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1581 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1584 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1594 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1600 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1607 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_1619 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1623 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1657 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_1669 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2893 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2905 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2911 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3341 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1147 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1161 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1185 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1197 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1203 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1241 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1253 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1259 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1273 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1297 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1353 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1365 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1371 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1377 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1416 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1429 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1441 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1448 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1460 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1470 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1480 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1505 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1508 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1518 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_1530 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_1538 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1553 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1571 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1583 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1615 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1627 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1639 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2827 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1007 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1021 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1045 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_105 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1057 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1063 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1077 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1101 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1119 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1213 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1225 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1263 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1275 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1287 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1299 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1311 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1319 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1323 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1331 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1336 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1353 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1382 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1394 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1398 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1412 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1422 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1432 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1442 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1454 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1461 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1473 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1501 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1509 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1513 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1517 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1539 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1551 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1555 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_1565 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1577 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_1589 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1603 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_1615 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2769 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2781 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2793 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2799 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2813 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2825 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2857 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2869 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2881 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2893 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2907 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2911 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_2921 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2927 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_2930 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2943 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2955 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3341 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1017 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1029 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1049 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1073 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1085 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1091 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1105 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1129 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1141 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1146 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1149 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1160 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1168 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1171 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1184 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1196 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1217 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1221 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1233 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1241 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1245 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1261 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1272 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1282 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1295 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1308 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1317 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1332 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1357 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1369 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1383 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1395 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1404 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1414 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_1426 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1429 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_1437 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1442 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1452 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1464 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_1476 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1489 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1492 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1502 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1514 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_1526 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1530 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2715 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2717 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2729 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2741 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2753 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2765 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2771 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2773 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2785 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2797 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2809 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2821 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2827 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2829 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2841 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2847 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2850 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2875 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2881 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_289 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2890 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2903 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_2916 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2920 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_2930 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_2938 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_973 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_979 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_993 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1001 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1007 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1015 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1027 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_1035 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1040 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1052 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1062 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1065 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1076 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1082 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1085 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1098 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1102 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1105 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1118 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1121 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1125 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1132 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1145 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1158 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1164 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1177 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1183 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1196 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1204 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1217 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1230 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1261 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1265 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1268 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1287 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1295 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1305 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1318 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1326 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1329 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1342 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_1345 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1356 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1366 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1379 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_1392 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1401 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_1413 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1420 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1432 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1444 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2701 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2713 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2725 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_273 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2737 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2743 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2745 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2757 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2769 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2773 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2776 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2784 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2789 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_2797 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2801 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2805 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2815 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2821 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2824 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2850 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2857 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2863 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_2876 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2880 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2890 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_2902 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_2910 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2913 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2937 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2949 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_2961 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3341 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_989 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1011 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1024 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1037 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1049 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1059 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1072 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1090 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1093 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1108 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1134 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1146 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1149 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1157 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1170 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1178 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1182 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1195 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1199 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1202 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1216 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1231 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1244 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1258 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1272 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1284 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_1292 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_1296 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_1304 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1309 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1315 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1329 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_1341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1347 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1359 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1371 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1385 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1421 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1427 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1465 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1477 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1483 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1497 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1521 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1533 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1539 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1553 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1577 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1589 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1595 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1609 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1633 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1651 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1665 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1701 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1707 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1721 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1745 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1757 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1763 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1765 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1777 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1801 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1813 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1819 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1821 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1833 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1857 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1869 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1875 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1877 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1889 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1913 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1925 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1931 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1933 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1945 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1969 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_1981 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_1987 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_1989 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2001 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2025 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2037 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2043 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2045 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2057 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2081 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2093 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2099 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2101 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2113 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2137 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2149 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2155 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2157 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2169 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2211 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2213 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2225 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2261 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2267 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2269 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2281 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2305 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2317 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2323 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2337 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2361 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2373 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2379 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2381 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2393 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2417 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2429 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2435 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2437 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2449 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2473 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2485 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2491 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2493 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2505 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2541 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2547 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2549 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2561 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2573 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2585 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2597 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2603 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2605 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2617 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2629 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_265 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2653 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2659 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2661 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2673 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2685 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2697 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2709 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2715 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2717 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2728 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2734 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2746 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2750 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2754 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_2770 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_2773 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2785 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2798 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2811 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_2824 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2829 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2841 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2853 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2865 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2877 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2883 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2885 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2897 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2909 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2921 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2933 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2939 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2953 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2965 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2977 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_2989 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_2995 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_2997 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3009 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3021 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3033 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3045 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3051 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3053 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3065 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3077 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3089 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3101 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3107 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3109 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3121 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3133 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3145 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3157 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3163 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3165 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3177 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3189 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3201 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3213 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3219 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3221 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3233 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3245 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3257 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3269 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3275 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3277 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3289 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3301 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3313 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3325 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3331 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3333 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3345 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3357 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3369 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3381 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3387 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3389 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3413 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3425 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3437 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3443 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3469 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3481 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3493 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3499 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3501 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3513 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3537 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3549 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3555 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3557 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3569 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3581 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3593 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3605 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3611 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3625 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3637 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3649 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3661 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3667 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3681 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3693 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3705 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3717 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3723 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3737 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3749 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3761 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3773 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3779 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3793 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3805 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3817 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3829 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3835 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3861 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3873 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3885 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3891 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3905 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3917 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3929 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3941 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_3947 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3973 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3985 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_3997 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4003 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4017 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4029 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4041 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4053 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4059 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4061 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4073 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4085 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4097 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4109 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4115 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4117 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4129 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4141 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4153 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4165 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4171 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4173 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4185 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4197 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4209 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4221 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4227 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4229 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4241 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4253 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4265 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4277 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4283 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4285 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4297 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4309 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4321 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4333 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4339 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4341 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4353 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4365 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4377 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4389 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4395 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4397 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4409 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4421 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4433 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4445 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4451 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4453 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4465 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4477 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4507 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4509 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4521 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4533 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4545 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4563 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4577 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4601 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4613 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4619 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4621 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4633 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4657 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4669 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4675 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4677 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4689 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_469 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4713 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4725 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4731 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4733 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4745 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4769 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4781 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4787 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4789 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4801 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4825 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4837 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4843 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4845 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4857 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4893 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4899 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4901 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4913 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4937 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_4949 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_4955 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4957 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4969 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4981 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_4993 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5005 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5011 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5013 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5025 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5037 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5049 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5061 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5067 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5069 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5081 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5093 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5105 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5117 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5123 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5125 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5137 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5149 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5161 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5173 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5179 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5181 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5193 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5205 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5217 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5229 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5235 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5237 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5249 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5261 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5273 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5285 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5291 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5293 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5305 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5317 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5329 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5341 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5347 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5349 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5361 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5373 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5385 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5397 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5403 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5405 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5417 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5429 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5441 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5453 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5459 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5461 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5473 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5485 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5497 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5509 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5515 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5517 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5529 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5541 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5553 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5565 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5571 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5573 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5585 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5597 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5609 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5621 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5627 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5629 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5641 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5653 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5665 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_5677 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_5683 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5685 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5697 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5709 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_5721 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_793 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_805 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_811 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_825 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_849 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_861 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_867 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_881 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_905 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_917 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_923 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_937 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_961 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_973 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_978 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_981 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_992 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_998 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1006 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_1009 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1021 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1034 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1047 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_105 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1060 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1065 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1071 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_1084 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1097 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1109 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1112 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1133 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1157 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1169 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1175 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1189 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1201 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1213 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1219 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_1222 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_1230 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1245 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1269 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1281 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1287 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1301 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1325 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1337 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1343 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1357 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1381 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1393 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1399 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1413 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1437 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1449 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1455 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1469 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1493 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1505 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1511 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1525 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1549 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1561 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1567 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1581 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1605 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1617 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1623 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1637 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1661 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1673 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1679 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1717 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1729 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1735 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1737 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1749 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1773 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1785 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1791 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1793 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1805 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1829 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1841 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1847 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1849 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1861 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1885 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1897 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1903 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1905 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1917 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1941 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_1953 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_1959 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1961 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1973 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_1997 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2009 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2015 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2017 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2029 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2053 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2065 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2071 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2073 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2085 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2097 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2109 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2121 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2127 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2129 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2141 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2165 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2177 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2183 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2185 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2197 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2209 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2221 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2233 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2239 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2241 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2253 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2277 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2289 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2295 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2297 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2309 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2333 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2345 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2351 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2353 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2365 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2389 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2401 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2407 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2409 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2421 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2445 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2457 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2463 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2465 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2477 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2489 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2501 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2513 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2519 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2521 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2533 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2557 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2569 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2575 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2577 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2589 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2613 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2625 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2631 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2633 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2645 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2657 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2669 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2681 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2687 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2689 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2703 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2716 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2729 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_273 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_2742 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2745 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2749 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2759 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2776 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2782 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2794 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2801 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2813 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2821 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2831 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2837 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2849 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2855 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2857 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2869 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2886 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2892 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2904 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2913 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_2925 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2931 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_2941 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2947 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_2959 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_2967 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2969 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2981 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_2993 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3005 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3017 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3023 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3025 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3037 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3049 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3061 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3073 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3079 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3081 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3093 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3105 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3117 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3129 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3135 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3137 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3149 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3161 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3173 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3185 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3191 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3193 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3205 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3217 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3229 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3241 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3247 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3249 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3261 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3273 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3285 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_329 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3297 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3303 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3305 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3317 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3329 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3341 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3353 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3359 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3373 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3385 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3397 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3409 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3415 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3441 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3453 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3465 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3471 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3497 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3509 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3521 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3527 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3553 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3565 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3577 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3583 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3597 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3609 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3621 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3633 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3639 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3653 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3665 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3677 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3689 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3695 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3709 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3721 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3733 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3745 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3751 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3765 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3777 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3789 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3801 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3807 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3821 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3833 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3845 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3857 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3863 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3877 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3889 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3901 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3913 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3919 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3933 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3945 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3957 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_3969 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_3975 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3977 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3989 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4001 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4013 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4025 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4031 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4033 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4045 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4057 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4069 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4081 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4087 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4089 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4101 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4113 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4125 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4137 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4143 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4145 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4157 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4169 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4181 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4193 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4199 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4201 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4213 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4225 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4237 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4249 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4255 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4257 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4269 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4281 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4293 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4305 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4311 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4313 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4325 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4337 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4349 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4361 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4367 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4369 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4381 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4393 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4405 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_441 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4417 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4423 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4425 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4437 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4461 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4473 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4479 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4481 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4493 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4517 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4529 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4535 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4537 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4549 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4573 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4585 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4591 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4593 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4605 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4629 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4641 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4647 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4649 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4661 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4685 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4697 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4703 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4705 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4717 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4741 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4753 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4759 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4761 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4773 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4797 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4809 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4815 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4817 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4829 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4853 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4865 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4871 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4873 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4885 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4909 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4921 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4927 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4929 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4941 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4953 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4965 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_497 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_4977 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_4983 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4985 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_4997 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5009 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5021 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5033 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5039 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5041 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5053 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5065 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5077 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5089 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5095 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5097 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5109 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5121 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5133 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5145 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5151 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5153 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5165 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5177 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5189 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5201 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5207 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5209 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5221 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5233 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5245 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5257 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5263 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5265 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5277 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5289 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5301 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5313 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5319 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5321 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5333 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5345 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5357 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5369 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5375 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5377 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5389 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5401 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5413 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5425 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5431 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5433 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5445 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5457 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5469 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5481 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5487 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5489 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5501 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5513 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5525 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5537 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5543 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5545 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5557 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5569 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5581 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5593 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5599 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5601 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5613 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5625 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5637 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5649 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5655 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5657 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5669 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5681 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5693 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_5705 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_5711 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_5713 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_5725 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_765 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_777 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_783 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_797 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_809 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_821 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_833 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_839 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_853 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_877 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_889 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_895 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_909 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_933 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_945 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_951 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_953 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_965 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_971 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_974 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_987 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_993 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_28 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_29 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_30 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_31 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_32 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_33 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_34 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_35 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_36 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_37 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_38 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_39 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_40 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_41 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_42 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_43 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_44 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_45 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_46 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_47 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_48 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_49 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_50 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_51 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_52 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_53 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_54 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_55 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_56 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_57 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_58 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_59 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_60 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_61 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_62 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_63 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_64 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_65 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_66 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_67 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_68 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_69 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_70 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_71 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_72 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_73 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_74 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_75 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_76 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__clkbuf_4 \u_rp[0].u_buf  (.A(ch_in[0]),
    .X(net91));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[100].u_buf  (.A(ch_in[100]),
    .X(net90));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[101].u_buf  (.A(ch_in[101]),
    .X(net89));
 sky130_fd_sc_hd__buf_2 \u_rp[102].u_buf  (.A(net161),
    .X(ch_out[102]));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[103].u_buf  (.A(ch_in[103]),
    .X(net88));
 sky130_fd_sc_hd__clkbuf_1 \u_rp[104].u_buf  (.A(ch_in[104]),
    .X(net87));
 sky130_fd_sc_hd__buf_2 \u_rp[105].u_buf  (.A(net160),
    .X(ch_out[105]));
 sky130_fd_sc_hd__buf_4 \u_rp[106].u_buf  (.A(ch_in[106]),
    .X(net86));
 sky130_fd_sc_hd__buf_2 \u_rp[107].u_buf  (.A(net159),
    .X(ch_out[107]));
 sky130_fd_sc_hd__buf_4 \u_rp[108].u_buf  (.A(ch_in[108]),
    .X(net85));
 sky130_fd_sc_hd__buf_2 \u_rp[109].u_buf  (.A(net158),
    .X(ch_out[109]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[10].u_buf  (.A(ch_in[10]),
    .X(net84));
 sky130_fd_sc_hd__buf_4 \u_rp[110].u_buf  (.A(ch_in[110]),
    .X(net83));
 sky130_fd_sc_hd__buf_2 \u_rp[111].u_buf  (.A(net157),
    .X(ch_out[111]));
 sky130_fd_sc_hd__buf_4 \u_rp[112].u_buf  (.A(ch_in[112]),
    .X(net82));
 sky130_fd_sc_hd__buf_2 \u_rp[113].u_buf  (.A(net156),
    .X(ch_out[113]));
 sky130_fd_sc_hd__buf_4 \u_rp[114].u_buf  (.A(ch_in[114]),
    .X(net81));
 sky130_fd_sc_hd__buf_2 \u_rp[115].u_buf  (.A(net155),
    .X(ch_out[115]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[116].u_buf  (.A(ch_in[116]),
    .X(net80));
 sky130_fd_sc_hd__buf_2 \u_rp[117].u_buf  (.A(net154),
    .X(ch_out[117]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[118].u_buf  (.A(ch_in[118]),
    .X(net79));
 sky130_fd_sc_hd__buf_2 \u_rp[119].u_buf  (.A(net153),
    .X(ch_out[119]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[11].u_buf  (.A(ch_in[11]),
    .X(net78));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[120].u_buf  (.A(ch_in[120]),
    .X(net77));
 sky130_fd_sc_hd__buf_2 \u_rp[121].u_buf  (.A(net152),
    .X(ch_out[121]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[122].u_buf  (.A(ch_in[122]),
    .X(net76));
 sky130_fd_sc_hd__buf_2 \u_rp[123].u_buf  (.A(net151),
    .X(ch_out[123]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[124].u_buf  (.A(ch_in[124]),
    .X(net75));
 sky130_fd_sc_hd__buf_2 \u_rp[125].u_buf  (.A(net150),
    .X(ch_out[125]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[126].u_buf  (.A(ch_in[126]),
    .X(net74));
 sky130_fd_sc_hd__buf_2 \u_rp[127].u_buf  (.A(net149),
    .X(ch_out[127]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[128].u_buf  (.A(ch_in[128]),
    .X(net73));
 sky130_fd_sc_hd__buf_2 \u_rp[129].u_buf  (.A(net148),
    .X(ch_out[129]));
 sky130_fd_sc_hd__buf_2 \u_rp[12].u_buf  (.A(net147),
    .X(ch_out[12]));
 sky130_fd_sc_hd__buf_2 \u_rp[130].u_buf  (.A(ch_in[130]),
    .X(net72));
 sky130_fd_sc_hd__buf_2 \u_rp[131].u_buf  (.A(net146),
    .X(ch_out[131]));
 sky130_fd_sc_hd__buf_2 \u_rp[132].u_buf  (.A(ch_in[132]),
    .X(net71));
 sky130_fd_sc_hd__buf_2 \u_rp[133].u_buf  (.A(net145),
    .X(ch_out[133]));
 sky130_fd_sc_hd__buf_2 \u_rp[134].u_buf  (.A(ch_in[134]),
    .X(net70));
 sky130_fd_sc_hd__buf_2 \u_rp[135].u_buf  (.A(net144),
    .X(ch_out[135]));
 sky130_fd_sc_hd__buf_2 \u_rp[136].u_buf  (.A(ch_in[136]),
    .X(net69));
 sky130_fd_sc_hd__buf_2 \u_rp[137].u_buf  (.A(net143),
    .X(ch_out[137]));
 sky130_fd_sc_hd__buf_2 \u_rp[138].u_buf  (.A(ch_in[138]),
    .X(net68));
 sky130_fd_sc_hd__buf_2 \u_rp[139].u_buf  (.A(net142),
    .X(ch_out[139]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[13].u_buf  (.A(ch_in[13]),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[140].u_buf  (.A(ch_in[140]),
    .X(net66));
 sky130_fd_sc_hd__buf_2 \u_rp[141].u_buf  (.A(net141),
    .X(ch_out[141]));
 sky130_fd_sc_hd__buf_2 \u_rp[142].u_buf  (.A(net140),
    .X(ch_out[142]));
 sky130_fd_sc_hd__buf_2 \u_rp[143].u_buf  (.A(net139),
    .X(ch_out[143]));
 sky130_fd_sc_hd__buf_2 \u_rp[144].u_buf  (.A(net138),
    .X(ch_out[144]));
 sky130_fd_sc_hd__buf_2 \u_rp[145].u_buf  (.A(net137),
    .X(ch_out[145]));
 sky130_fd_sc_hd__buf_2 \u_rp[146].u_buf  (.A(net136),
    .X(ch_out[146]));
 sky130_fd_sc_hd__buf_2 \u_rp[147].u_buf  (.A(net135),
    .X(ch_out[147]));
 sky130_fd_sc_hd__buf_2 \u_rp[148].u_buf  (.A(net134),
    .X(ch_out[148]));
 sky130_fd_sc_hd__buf_2 \u_rp[149].u_buf  (.A(net133),
    .X(ch_out[149]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[14].u_buf  (.A(ch_in[14]),
    .X(net65));
 sky130_fd_sc_hd__buf_2 \u_rp[150].u_buf  (.A(net132),
    .X(ch_out[150]));
 sky130_fd_sc_hd__buf_2 \u_rp[151].u_buf  (.A(net131),
    .X(ch_out[151]));
 sky130_fd_sc_hd__buf_2 \u_rp[152].u_buf  (.A(net130),
    .X(ch_out[152]));
 sky130_fd_sc_hd__buf_2 \u_rp[153].u_buf  (.A(net129),
    .X(ch_out[153]));
 sky130_fd_sc_hd__buf_2 \u_rp[154].u_buf  (.A(net128),
    .X(ch_out[154]));
 sky130_fd_sc_hd__buf_2 \u_rp[155].u_buf  (.A(net127),
    .X(ch_out[155]));
 sky130_fd_sc_hd__buf_2 \u_rp[156].u_buf  (.A(net126),
    .X(ch_out[156]));
 sky130_fd_sc_hd__buf_2 \u_rp[157].u_buf  (.A(net125),
    .X(ch_out[157]));
 sky130_fd_sc_hd__buf_2 \u_rp[158].u_buf  (.A(net124),
    .X(ch_out[158]));
 sky130_fd_sc_hd__buf_2 \u_rp[159].u_buf  (.A(net123),
    .X(ch_out[159]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[15].u_buf  (.A(ch_in[15]),
    .X(net64));
 sky130_fd_sc_hd__buf_2 \u_rp[160].u_buf  (.A(net122),
    .X(ch_out[160]));
 sky130_fd_sc_hd__buf_2 \u_rp[161].u_buf  (.A(ch_in[161]),
    .X(ch_out[161]));
 sky130_fd_sc_hd__buf_2 \u_rp[162].u_buf  (.A(ch_in[162]),
    .X(ch_out[162]));
 sky130_fd_sc_hd__buf_2 \u_rp[163].u_buf  (.A(ch_in[163]),
    .X(ch_out[163]));
 sky130_fd_sc_hd__buf_2 \u_rp[164].u_buf  (.A(ch_in[164]),
    .X(ch_out[164]));
 sky130_fd_sc_hd__buf_2 \u_rp[165].u_buf  (.A(ch_in[165]),
    .X(ch_out[165]));
 sky130_fd_sc_hd__buf_2 \u_rp[166].u_buf  (.A(ch_in[166]),
    .X(ch_out[166]));
 sky130_fd_sc_hd__buf_2 \u_rp[167].u_buf  (.A(ch_in[167]),
    .X(ch_out[167]));
 sky130_fd_sc_hd__buf_2 \u_rp[168].u_buf  (.A(ch_in[168]),
    .X(ch_out[168]));
 sky130_fd_sc_hd__buf_2 \u_rp[169].u_buf  (.A(ch_in[169]),
    .X(ch_out[169]));
 sky130_fd_sc_hd__buf_2 \u_rp[16].u_buf  (.A(net121),
    .X(ch_out[16]));
 sky130_fd_sc_hd__buf_2 \u_rp[170].u_buf  (.A(ch_in[170]),
    .X(ch_out[170]));
 sky130_fd_sc_hd__buf_2 \u_rp[171].u_buf  (.A(ch_in[171]),
    .X(ch_out[171]));
 sky130_fd_sc_hd__buf_2 \u_rp[172].u_buf  (.A(ch_in[172]),
    .X(ch_out[172]));
 sky130_fd_sc_hd__buf_2 \u_rp[173].u_buf  (.A(ch_in[173]),
    .X(ch_out[173]));
 sky130_fd_sc_hd__buf_2 \u_rp[174].u_buf  (.A(ch_in[174]),
    .X(ch_out[174]));
 sky130_fd_sc_hd__buf_2 \u_rp[175].u_buf  (.A(ch_in[175]),
    .X(ch_out[175]));
 sky130_fd_sc_hd__buf_2 \u_rp[176].u_buf  (.A(ch_in[176]),
    .X(ch_out[176]));
 sky130_fd_sc_hd__buf_2 \u_rp[177].u_buf  (.A(ch_in[177]),
    .X(ch_out[177]));
 sky130_fd_sc_hd__buf_2 \u_rp[178].u_buf  (.A(ch_in[178]),
    .X(ch_out[178]));
 sky130_fd_sc_hd__buf_2 \u_rp[179].u_buf  (.A(ch_in[179]),
    .X(ch_out[179]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[17].u_buf  (.A(ch_in[17]),
    .X(net63));
 sky130_fd_sc_hd__buf_2 \u_rp[180].u_buf  (.A(ch_in[180]),
    .X(ch_out[180]));
 sky130_fd_sc_hd__buf_2 \u_rp[181].u_buf  (.A(ch_in[181]),
    .X(ch_out[181]));
 sky130_fd_sc_hd__buf_2 \u_rp[182].u_buf  (.A(ch_in[182]),
    .X(ch_out[182]));
 sky130_fd_sc_hd__buf_2 \u_rp[183].u_buf  (.A(ch_in[183]),
    .X(ch_out[183]));
 sky130_fd_sc_hd__buf_2 \u_rp[184].u_buf  (.A(ch_in[184]),
    .X(ch_out[184]));
 sky130_fd_sc_hd__buf_2 \u_rp[185].u_buf  (.A(ch_in[185]),
    .X(ch_out[185]));
 sky130_fd_sc_hd__buf_2 \u_rp[186].u_buf  (.A(ch_in[186]),
    .X(ch_out[186]));
 sky130_fd_sc_hd__buf_2 \u_rp[187].u_buf  (.A(ch_in[187]),
    .X(ch_out[187]));
 sky130_fd_sc_hd__buf_2 \u_rp[188].u_buf  (.A(ch_in[188]),
    .X(ch_out[188]));
 sky130_fd_sc_hd__buf_2 \u_rp[189].u_buf  (.A(ch_in[189]),
    .X(ch_out[189]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[18].u_buf  (.A(ch_in[18]),
    .X(net62));
 sky130_fd_sc_hd__buf_2 \u_rp[190].u_buf  (.A(ch_in[190]),
    .X(ch_out[190]));
 sky130_fd_sc_hd__buf_2 \u_rp[191].u_buf  (.A(ch_in[191]),
    .X(ch_out[191]));
 sky130_fd_sc_hd__buf_2 \u_rp[192].u_buf  (.A(ch_in[192]),
    .X(ch_out[192]));
 sky130_fd_sc_hd__buf_2 \u_rp[193].u_buf  (.A(ch_in[193]),
    .X(ch_out[193]));
 sky130_fd_sc_hd__buf_2 \u_rp[194].u_buf  (.A(ch_in[194]),
    .X(ch_out[194]));
 sky130_fd_sc_hd__buf_2 \u_rp[195].u_buf  (.A(ch_in[195]),
    .X(ch_out[195]));
 sky130_fd_sc_hd__buf_2 \u_rp[196].u_buf  (.A(ch_in[196]),
    .X(ch_out[196]));
 sky130_fd_sc_hd__buf_2 \u_rp[197].u_buf  (.A(ch_in[197]),
    .X(ch_out[197]));
 sky130_fd_sc_hd__buf_2 \u_rp[198].u_buf  (.A(ch_in[198]),
    .X(ch_out[198]));
 sky130_fd_sc_hd__buf_2 \u_rp[199].u_buf  (.A(ch_in[199]),
    .X(ch_out[199]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[19].u_buf  (.A(ch_in[19]),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[1].u_buf  (.A(ch_in[1]),
    .X(net60));
 sky130_fd_sc_hd__buf_2 \u_rp[200].u_buf  (.A(ch_in[200]),
    .X(ch_out[200]));
 sky130_fd_sc_hd__buf_2 \u_rp[201].u_buf  (.A(ch_in[201]),
    .X(ch_out[201]));
 sky130_fd_sc_hd__buf_2 \u_rp[202].u_buf  (.A(ch_in[202]),
    .X(ch_out[202]));
 sky130_fd_sc_hd__buf_2 \u_rp[203].u_buf  (.A(ch_in[203]),
    .X(ch_out[203]));
 sky130_fd_sc_hd__buf_2 \u_rp[204].u_buf  (.A(ch_in[204]),
    .X(ch_out[204]));
 sky130_fd_sc_hd__buf_2 \u_rp[205].u_buf  (.A(ch_in[205]),
    .X(ch_out[205]));
 sky130_fd_sc_hd__buf_2 \u_rp[206].u_buf  (.A(ch_in[206]),
    .X(ch_out[206]));
 sky130_fd_sc_hd__buf_2 \u_rp[207].u_buf  (.A(ch_in[207]),
    .X(ch_out[207]));
 sky130_fd_sc_hd__buf_2 \u_rp[208].u_buf  (.A(ch_in[208]),
    .X(ch_out[208]));
 sky130_fd_sc_hd__buf_2 \u_rp[209].u_buf  (.A(ch_in[209]),
    .X(ch_out[209]));
 sky130_fd_sc_hd__buf_2 \u_rp[20].u_buf  (.A(net120),
    .X(ch_out[20]));
 sky130_fd_sc_hd__buf_2 \u_rp[210].u_buf  (.A(ch_in[210]),
    .X(ch_out[210]));
 sky130_fd_sc_hd__buf_2 \u_rp[211].u_buf  (.A(ch_in[211]),
    .X(ch_out[211]));
 sky130_fd_sc_hd__buf_2 \u_rp[212].u_buf  (.A(ch_in[212]),
    .X(ch_out[212]));
 sky130_fd_sc_hd__buf_2 \u_rp[213].u_buf  (.A(ch_in[213]),
    .X(ch_out[213]));
 sky130_fd_sc_hd__buf_2 \u_rp[214].u_buf  (.A(ch_in[214]),
    .X(ch_out[214]));
 sky130_fd_sc_hd__buf_2 \u_rp[215].u_buf  (.A(ch_in[215]),
    .X(ch_out[215]));
 sky130_fd_sc_hd__buf_2 \u_rp[216].u_buf  (.A(ch_in[216]),
    .X(ch_out[216]));
 sky130_fd_sc_hd__buf_2 \u_rp[217].u_buf  (.A(ch_in[217]),
    .X(ch_out[217]));
 sky130_fd_sc_hd__buf_2 \u_rp[218].u_buf  (.A(ch_in[218]),
    .X(ch_out[218]));
 sky130_fd_sc_hd__buf_2 \u_rp[219].u_buf  (.A(ch_in[219]),
    .X(ch_out[219]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[21].u_buf  (.A(ch_in[21]),
    .X(net59));
 sky130_fd_sc_hd__buf_2 \u_rp[220].u_buf  (.A(ch_in[220]),
    .X(ch_out[220]));
 sky130_fd_sc_hd__buf_2 \u_rp[221].u_buf  (.A(ch_in[221]),
    .X(ch_out[221]));
 sky130_fd_sc_hd__buf_2 \u_rp[222].u_buf  (.A(ch_in[222]),
    .X(ch_out[222]));
 sky130_fd_sc_hd__buf_2 \u_rp[223].u_buf  (.A(ch_in[223]),
    .X(ch_out[223]));
 sky130_fd_sc_hd__buf_2 \u_rp[224].u_buf  (.A(ch_in[224]),
    .X(ch_out[224]));
 sky130_fd_sc_hd__buf_2 \u_rp[225].u_buf  (.A(ch_in[225]),
    .X(ch_out[225]));
 sky130_fd_sc_hd__buf_2 \u_rp[226].u_buf  (.A(ch_in[226]),
    .X(ch_out[226]));
 sky130_fd_sc_hd__buf_2 \u_rp[227].u_buf  (.A(ch_in[227]),
    .X(ch_out[227]));
 sky130_fd_sc_hd__buf_2 \u_rp[228].u_buf  (.A(ch_in[228]),
    .X(ch_out[228]));
 sky130_fd_sc_hd__buf_2 \u_rp[229].u_buf  (.A(ch_in[229]),
    .X(ch_out[229]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[22].u_buf  (.A(ch_in[22]),
    .X(net58));
 sky130_fd_sc_hd__buf_2 \u_rp[230].u_buf  (.A(ch_in[230]),
    .X(ch_out[230]));
 sky130_fd_sc_hd__buf_2 \u_rp[231].u_buf  (.A(ch_in[231]),
    .X(ch_out[231]));
 sky130_fd_sc_hd__buf_2 \u_rp[232].u_buf  (.A(ch_in[232]),
    .X(ch_out[232]));
 sky130_fd_sc_hd__buf_2 \u_rp[233].u_buf  (.A(ch_in[233]),
    .X(ch_out[233]));
 sky130_fd_sc_hd__buf_2 \u_rp[234].u_buf  (.A(ch_in[234]),
    .X(ch_out[234]));
 sky130_fd_sc_hd__buf_2 \u_rp[235].u_buf  (.A(ch_in[235]),
    .X(ch_out[235]));
 sky130_fd_sc_hd__buf_2 \u_rp[236].u_buf  (.A(ch_in[236]),
    .X(ch_out[236]));
 sky130_fd_sc_hd__buf_2 \u_rp[237].u_buf  (.A(ch_in[237]),
    .X(ch_out[237]));
 sky130_fd_sc_hd__buf_2 \u_rp[238].u_buf  (.A(ch_in[238]),
    .X(ch_out[238]));
 sky130_fd_sc_hd__buf_2 \u_rp[239].u_buf  (.A(ch_in[239]),
    .X(ch_out[239]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[23].u_buf  (.A(ch_in[23]),
    .X(net57));
 sky130_fd_sc_hd__buf_2 \u_rp[240].u_buf  (.A(ch_in[240]),
    .X(ch_out[240]));
 sky130_fd_sc_hd__buf_2 \u_rp[241].u_buf  (.A(ch_in[241]),
    .X(ch_out[241]));
 sky130_fd_sc_hd__buf_2 \u_rp[242].u_buf  (.A(ch_in[242]),
    .X(ch_out[242]));
 sky130_fd_sc_hd__buf_2 \u_rp[243].u_buf  (.A(ch_in[243]),
    .X(ch_out[243]));
 sky130_fd_sc_hd__buf_2 \u_rp[244].u_buf  (.A(ch_in[244]),
    .X(ch_out[244]));
 sky130_fd_sc_hd__buf_2 \u_rp[245].u_buf  (.A(ch_in[245]),
    .X(ch_out[245]));
 sky130_fd_sc_hd__buf_2 \u_rp[246].u_buf  (.A(ch_in[246]),
    .X(ch_out[246]));
 sky130_fd_sc_hd__buf_2 \u_rp[247].u_buf  (.A(ch_in[247]),
    .X(ch_out[247]));
 sky130_fd_sc_hd__buf_2 \u_rp[248].u_buf  (.A(ch_in[248]),
    .X(ch_out[248]));
 sky130_fd_sc_hd__buf_2 \u_rp[249].u_buf  (.A(ch_in[249]),
    .X(ch_out[249]));
 sky130_fd_sc_hd__buf_2 \u_rp[24].u_buf  (.A(net119),
    .X(ch_out[24]));
 sky130_fd_sc_hd__buf_2 \u_rp[250].u_buf  (.A(ch_in[250]),
    .X(ch_out[250]));
 sky130_fd_sc_hd__buf_2 \u_rp[251].u_buf  (.A(ch_in[251]),
    .X(ch_out[251]));
 sky130_fd_sc_hd__buf_2 \u_rp[252].u_buf  (.A(ch_in[252]),
    .X(ch_out[252]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[25].u_buf  (.A(ch_in[25]),
    .X(net56));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[26].u_buf  (.A(ch_in[26]),
    .X(net55));
 sky130_fd_sc_hd__buf_2 \u_rp[27].u_buf  (.A(net118),
    .X(ch_out[27]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[28].u_buf  (.A(ch_in[28]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[29].u_buf  (.A(ch_in[29]),
    .X(net53));
 sky130_fd_sc_hd__buf_2 \u_rp[2].u_buf  (.A(net117),
    .X(ch_out[2]));
 sky130_fd_sc_hd__buf_2 \u_rp[30].u_buf  (.A(net116),
    .X(ch_out[30]));
 sky130_fd_sc_hd__buf_2 \u_rp[31].u_buf  (.A(ch_in[31]),
    .X(net52));
 sky130_fd_sc_hd__buf_2 \u_rp[32].u_buf  (.A(ch_in[32]),
    .X(net51));
 sky130_fd_sc_hd__buf_2 \u_rp[33].u_buf  (.A(net115),
    .X(ch_out[33]));
 sky130_fd_sc_hd__buf_2 \u_rp[34].u_buf  (.A(ch_in[34]),
    .X(net50));
 sky130_fd_sc_hd__buf_2 \u_rp[35].u_buf  (.A(ch_in[35]),
    .X(net49));
 sky130_fd_sc_hd__buf_2 \u_rp[36].u_buf  (.A(net114),
    .X(ch_out[36]));
 sky130_fd_sc_hd__buf_2 \u_rp[37].u_buf  (.A(ch_in[37]),
    .X(net48));
 sky130_fd_sc_hd__buf_2 \u_rp[38].u_buf  (.A(ch_in[38]),
    .X(net47));
 sky130_fd_sc_hd__buf_2 \u_rp[39].u_buf  (.A(net113),
    .X(ch_out[39]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[3].u_buf  (.A(ch_in[3]),
    .X(net46));
 sky130_fd_sc_hd__buf_2 \u_rp[40].u_buf  (.A(ch_in[40]),
    .X(net45));
 sky130_fd_sc_hd__buf_2 \u_rp[41].u_buf  (.A(ch_in[41]),
    .X(net44));
 sky130_fd_sc_hd__buf_2 \u_rp[42].u_buf  (.A(net112),
    .X(ch_out[42]));
 sky130_fd_sc_hd__buf_2 \u_rp[43].u_buf  (.A(ch_in[43]),
    .X(net43));
 sky130_fd_sc_hd__buf_2 \u_rp[44].u_buf  (.A(ch_in[44]),
    .X(net42));
 sky130_fd_sc_hd__buf_2 \u_rp[45].u_buf  (.A(net111),
    .X(ch_out[45]));
 sky130_fd_sc_hd__buf_2 \u_rp[46].u_buf  (.A(ch_in[46]),
    .X(net41));
 sky130_fd_sc_hd__buf_2 \u_rp[47].u_buf  (.A(ch_in[47]),
    .X(net40));
 sky130_fd_sc_hd__buf_2 \u_rp[48].u_buf  (.A(net110),
    .X(ch_out[48]));
 sky130_fd_sc_hd__buf_2 \u_rp[49].u_buf  (.A(ch_in[49]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[4].u_buf  (.A(ch_in[4]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 \u_rp[50].u_buf  (.A(ch_in[50]),
    .X(net37));
 sky130_fd_sc_hd__buf_2 \u_rp[51].u_buf  (.A(net109),
    .X(ch_out[51]));
 sky130_fd_sc_hd__buf_2 \u_rp[52].u_buf  (.A(ch_in[52]),
    .X(net36));
 sky130_fd_sc_hd__buf_2 \u_rp[53].u_buf  (.A(ch_in[53]),
    .X(net35));
 sky130_fd_sc_hd__buf_2 \u_rp[54].u_buf  (.A(net108),
    .X(ch_out[54]));
 sky130_fd_sc_hd__buf_2 \u_rp[55].u_buf  (.A(ch_in[55]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 \u_rp[56].u_buf  (.A(ch_in[56]),
    .X(net33));
 sky130_fd_sc_hd__buf_2 \u_rp[57].u_buf  (.A(net107),
    .X(ch_out[57]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[58].u_buf  (.A(ch_in[58]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[59].u_buf  (.A(ch_in[59]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[5].u_buf  (.A(ch_in[5]),
    .X(net30));
 sky130_fd_sc_hd__buf_2 \u_rp[60].u_buf  (.A(net106),
    .X(ch_out[60]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[61].u_buf  (.A(ch_in[61]),
    .X(net29));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[62].u_buf  (.A(ch_in[62]),
    .X(net28));
 sky130_fd_sc_hd__buf_2 \u_rp[63].u_buf  (.A(net105),
    .X(ch_out[63]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[64].u_buf  (.A(ch_in[64]),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[65].u_buf  (.A(ch_in[65]),
    .X(net26));
 sky130_fd_sc_hd__buf_2 \u_rp[66].u_buf  (.A(net104),
    .X(ch_out[66]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[67].u_buf  (.A(ch_in[67]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[68].u_buf  (.A(ch_in[68]),
    .X(net24));
 sky130_fd_sc_hd__buf_2 \u_rp[69].u_buf  (.A(net103),
    .X(ch_out[69]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[6].u_buf  (.A(ch_in[6]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[70].u_buf  (.A(ch_in[70]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[71].u_buf  (.A(ch_in[71]),
    .X(net21));
 sky130_fd_sc_hd__buf_2 \u_rp[72].u_buf  (.A(net102),
    .X(ch_out[72]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[73].u_buf  (.A(ch_in[73]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[74].u_buf  (.A(ch_in[74]),
    .X(net19));
 sky130_fd_sc_hd__buf_2 \u_rp[75].u_buf  (.A(net101),
    .X(ch_out[75]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[76].u_buf  (.A(ch_in[76]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[77].u_buf  (.A(ch_in[77]),
    .X(net17));
 sky130_fd_sc_hd__buf_2 \u_rp[78].u_buf  (.A(net100),
    .X(ch_out[78]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[79].u_buf  (.A(ch_in[79]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[7].u_buf  (.A(ch_in[7]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[80].u_buf  (.A(ch_in[80]),
    .X(net14));
 sky130_fd_sc_hd__buf_2 \u_rp[81].u_buf  (.A(net99),
    .X(ch_out[81]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[82].u_buf  (.A(ch_in[82]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[83].u_buf  (.A(ch_in[83]),
    .X(net12));
 sky130_fd_sc_hd__buf_2 \u_rp[84].u_buf  (.A(net98),
    .X(ch_out[84]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[85].u_buf  (.A(ch_in[85]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[86].u_buf  (.A(ch_in[86]),
    .X(net10));
 sky130_fd_sc_hd__buf_2 \u_rp[87].u_buf  (.A(net97),
    .X(ch_out[87]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[88].u_buf  (.A(ch_in[88]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[89].u_buf  (.A(ch_in[89]),
    .X(net8));
 sky130_fd_sc_hd__buf_2 \u_rp[8].u_buf  (.A(net96),
    .X(ch_out[8]));
 sky130_fd_sc_hd__buf_2 \u_rp[90].u_buf  (.A(net95),
    .X(ch_out[90]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[91].u_buf  (.A(ch_in[91]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[92].u_buf  (.A(ch_in[92]),
    .X(net6));
 sky130_fd_sc_hd__buf_2 \u_rp[93].u_buf  (.A(net94),
    .X(ch_out[93]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[94].u_buf  (.A(ch_in[94]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[95].u_buf  (.A(ch_in[95]),
    .X(net4));
 sky130_fd_sc_hd__buf_2 \u_rp[96].u_buf  (.A(net93),
    .X(ch_out[96]));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[97].u_buf  (.A(ch_in[97]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 \u_rp[98].u_buf  (.A(ch_in[98]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 \u_rp[99].u_buf  (.A(net92),
    .X(ch_out[99]));
 sky130_fd_sc_hd__clkbuf_4 \u_rp[9].u_buf  (.A(ch_in[9]),
    .X(net1));
 sky130_fd_sc_hd__buf_6 wire1 (.A(net1),
    .X(ch_out[9]));
 sky130_fd_sc_hd__buf_4 wire10 (.A(net10),
    .X(ch_out[86]));
 sky130_fd_sc_hd__buf_4 wire100 (.A(ch_in[78]),
    .X(net100));
 sky130_fd_sc_hd__buf_4 wire101 (.A(ch_in[75]),
    .X(net101));
 sky130_fd_sc_hd__buf_6 wire102 (.A(ch_in[72]),
    .X(net102));
 sky130_fd_sc_hd__buf_6 wire103 (.A(ch_in[69]),
    .X(net103));
 sky130_fd_sc_hd__buf_6 wire104 (.A(ch_in[66]),
    .X(net104));
 sky130_fd_sc_hd__buf_6 wire105 (.A(ch_in[63]),
    .X(net105));
 sky130_fd_sc_hd__buf_6 wire106 (.A(ch_in[60]),
    .X(net106));
 sky130_fd_sc_hd__buf_6 wire107 (.A(ch_in[57]),
    .X(net107));
 sky130_fd_sc_hd__buf_6 wire108 (.A(ch_in[54]),
    .X(net108));
 sky130_fd_sc_hd__buf_6 wire109 (.A(ch_in[51]),
    .X(net109));
 sky130_fd_sc_hd__buf_4 wire11 (.A(net11),
    .X(ch_out[85]));
 sky130_fd_sc_hd__buf_6 wire110 (.A(ch_in[48]),
    .X(net110));
 sky130_fd_sc_hd__buf_6 wire111 (.A(ch_in[45]),
    .X(net111));
 sky130_fd_sc_hd__buf_6 wire112 (.A(ch_in[42]),
    .X(net112));
 sky130_fd_sc_hd__buf_6 wire113 (.A(ch_in[39]),
    .X(net113));
 sky130_fd_sc_hd__buf_6 wire114 (.A(ch_in[36]),
    .X(net114));
 sky130_fd_sc_hd__buf_6 wire115 (.A(ch_in[33]),
    .X(net115));
 sky130_fd_sc_hd__buf_6 wire116 (.A(ch_in[30]),
    .X(net116));
 sky130_fd_sc_hd__buf_6 wire117 (.A(ch_in[2]),
    .X(net117));
 sky130_fd_sc_hd__buf_6 wire118 (.A(ch_in[27]),
    .X(net118));
 sky130_fd_sc_hd__buf_6 wire119 (.A(ch_in[24]),
    .X(net119));
 sky130_fd_sc_hd__buf_4 wire12 (.A(net12),
    .X(ch_out[83]));
 sky130_fd_sc_hd__buf_6 wire120 (.A(ch_in[20]),
    .X(net120));
 sky130_fd_sc_hd__buf_6 wire121 (.A(ch_in[16]),
    .X(net121));
 sky130_fd_sc_hd__buf_4 wire122 (.A(ch_in[160]),
    .X(net122));
 sky130_fd_sc_hd__buf_4 wire123 (.A(ch_in[159]),
    .X(net123));
 sky130_fd_sc_hd__buf_4 wire124 (.A(ch_in[158]),
    .X(net124));
 sky130_fd_sc_hd__buf_4 wire125 (.A(ch_in[157]),
    .X(net125));
 sky130_fd_sc_hd__buf_4 wire126 (.A(ch_in[156]),
    .X(net126));
 sky130_fd_sc_hd__buf_4 wire127 (.A(ch_in[155]),
    .X(net127));
 sky130_fd_sc_hd__buf_4 wire128 (.A(ch_in[154]),
    .X(net128));
 sky130_fd_sc_hd__buf_4 wire129 (.A(ch_in[153]),
    .X(net129));
 sky130_fd_sc_hd__buf_4 wire13 (.A(net13),
    .X(ch_out[82]));
 sky130_fd_sc_hd__buf_4 wire130 (.A(ch_in[152]),
    .X(net130));
 sky130_fd_sc_hd__buf_4 wire131 (.A(ch_in[151]),
    .X(net131));
 sky130_fd_sc_hd__buf_4 wire132 (.A(ch_in[150]),
    .X(net132));
 sky130_fd_sc_hd__buf_4 wire133 (.A(ch_in[149]),
    .X(net133));
 sky130_fd_sc_hd__buf_4 wire134 (.A(ch_in[148]),
    .X(net134));
 sky130_fd_sc_hd__buf_4 wire135 (.A(ch_in[147]),
    .X(net135));
 sky130_fd_sc_hd__buf_4 wire136 (.A(ch_in[146]),
    .X(net136));
 sky130_fd_sc_hd__buf_4 wire137 (.A(ch_in[145]),
    .X(net137));
 sky130_fd_sc_hd__buf_6 wire138 (.A(ch_in[144]),
    .X(net138));
 sky130_fd_sc_hd__buf_6 wire139 (.A(ch_in[143]),
    .X(net139));
 sky130_fd_sc_hd__buf_4 wire14 (.A(net14),
    .X(ch_out[80]));
 sky130_fd_sc_hd__buf_6 wire140 (.A(ch_in[142]),
    .X(net140));
 sky130_fd_sc_hd__buf_6 wire141 (.A(ch_in[141]),
    .X(net141));
 sky130_fd_sc_hd__buf_6 wire142 (.A(ch_in[139]),
    .X(net142));
 sky130_fd_sc_hd__buf_6 wire143 (.A(ch_in[137]),
    .X(net143));
 sky130_fd_sc_hd__buf_6 wire144 (.A(ch_in[135]),
    .X(net144));
 sky130_fd_sc_hd__buf_6 wire145 (.A(ch_in[133]),
    .X(net145));
 sky130_fd_sc_hd__buf_6 wire146 (.A(ch_in[131]),
    .X(net146));
 sky130_fd_sc_hd__buf_6 wire147 (.A(ch_in[12]),
    .X(net147));
 sky130_fd_sc_hd__buf_6 wire148 (.A(ch_in[129]),
    .X(net148));
 sky130_fd_sc_hd__buf_6 wire149 (.A(ch_in[127]),
    .X(net149));
 sky130_fd_sc_hd__buf_6 wire15 (.A(net15),
    .X(ch_out[7]));
 sky130_fd_sc_hd__buf_6 wire150 (.A(ch_in[125]),
    .X(net150));
 sky130_fd_sc_hd__buf_6 wire151 (.A(ch_in[123]),
    .X(net151));
 sky130_fd_sc_hd__buf_6 wire152 (.A(ch_in[121]),
    .X(net152));
 sky130_fd_sc_hd__buf_6 wire153 (.A(ch_in[119]),
    .X(net153));
 sky130_fd_sc_hd__buf_6 wire154 (.A(ch_in[117]),
    .X(net154));
 sky130_fd_sc_hd__buf_6 wire155 (.A(ch_in[115]),
    .X(net155));
 sky130_fd_sc_hd__buf_6 wire156 (.A(ch_in[113]),
    .X(net156));
 sky130_fd_sc_hd__buf_6 wire157 (.A(ch_in[111]),
    .X(net157));
 sky130_fd_sc_hd__buf_6 wire158 (.A(ch_in[109]),
    .X(net158));
 sky130_fd_sc_hd__buf_6 wire159 (.A(ch_in[107]),
    .X(net159));
 sky130_fd_sc_hd__buf_4 wire16 (.A(net16),
    .X(ch_out[79]));
 sky130_fd_sc_hd__buf_4 wire160 (.A(ch_in[105]),
    .X(net160));
 sky130_fd_sc_hd__buf_4 wire161 (.A(ch_in[102]),
    .X(net161));
 sky130_fd_sc_hd__buf_4 wire17 (.A(net17),
    .X(ch_out[77]));
 sky130_fd_sc_hd__buf_4 wire18 (.A(net18),
    .X(ch_out[76]));
 sky130_fd_sc_hd__buf_4 wire19 (.A(net19),
    .X(ch_out[74]));
 sky130_fd_sc_hd__buf_4 wire2 (.A(net2),
    .X(ch_out[98]));
 sky130_fd_sc_hd__buf_4 wire20 (.A(net20),
    .X(ch_out[73]));
 sky130_fd_sc_hd__buf_4 wire21 (.A(net21),
    .X(ch_out[71]));
 sky130_fd_sc_hd__buf_4 wire22 (.A(net22),
    .X(ch_out[70]));
 sky130_fd_sc_hd__buf_6 wire23 (.A(net23),
    .X(ch_out[6]));
 sky130_fd_sc_hd__buf_6 wire24 (.A(net24),
    .X(ch_out[68]));
 sky130_fd_sc_hd__buf_6 wire25 (.A(net25),
    .X(ch_out[67]));
 sky130_fd_sc_hd__buf_6 wire26 (.A(net26),
    .X(ch_out[65]));
 sky130_fd_sc_hd__buf_6 wire27 (.A(net27),
    .X(ch_out[64]));
 sky130_fd_sc_hd__buf_6 wire28 (.A(net28),
    .X(ch_out[62]));
 sky130_fd_sc_hd__buf_6 wire29 (.A(net29),
    .X(ch_out[61]));
 sky130_fd_sc_hd__buf_4 wire3 (.A(net3),
    .X(ch_out[97]));
 sky130_fd_sc_hd__buf_6 wire30 (.A(net30),
    .X(ch_out[5]));
 sky130_fd_sc_hd__buf_6 wire31 (.A(net31),
    .X(ch_out[59]));
 sky130_fd_sc_hd__buf_6 wire32 (.A(net32),
    .X(ch_out[58]));
 sky130_fd_sc_hd__buf_6 wire33 (.A(net33),
    .X(ch_out[56]));
 sky130_fd_sc_hd__buf_6 wire34 (.A(net34),
    .X(ch_out[55]));
 sky130_fd_sc_hd__buf_6 wire35 (.A(net35),
    .X(ch_out[53]));
 sky130_fd_sc_hd__buf_6 wire36 (.A(net36),
    .X(ch_out[52]));
 sky130_fd_sc_hd__buf_6 wire37 (.A(net37),
    .X(ch_out[50]));
 sky130_fd_sc_hd__buf_6 wire38 (.A(net38),
    .X(ch_out[4]));
 sky130_fd_sc_hd__buf_6 wire39 (.A(net39),
    .X(ch_out[49]));
 sky130_fd_sc_hd__buf_4 wire4 (.A(net4),
    .X(ch_out[95]));
 sky130_fd_sc_hd__buf_6 wire40 (.A(net40),
    .X(ch_out[47]));
 sky130_fd_sc_hd__buf_6 wire41 (.A(net41),
    .X(ch_out[46]));
 sky130_fd_sc_hd__buf_6 wire42 (.A(net42),
    .X(ch_out[44]));
 sky130_fd_sc_hd__buf_6 wire43 (.A(net43),
    .X(ch_out[43]));
 sky130_fd_sc_hd__buf_6 wire44 (.A(net44),
    .X(ch_out[41]));
 sky130_fd_sc_hd__buf_6 wire45 (.A(net45),
    .X(ch_out[40]));
 sky130_fd_sc_hd__buf_6 wire46 (.A(net46),
    .X(ch_out[3]));
 sky130_fd_sc_hd__buf_6 wire47 (.A(net47),
    .X(ch_out[38]));
 sky130_fd_sc_hd__buf_6 wire48 (.A(net48),
    .X(ch_out[37]));
 sky130_fd_sc_hd__buf_6 wire49 (.A(net49),
    .X(ch_out[35]));
 sky130_fd_sc_hd__buf_4 wire5 (.A(net5),
    .X(ch_out[94]));
 sky130_fd_sc_hd__buf_6 wire50 (.A(net50),
    .X(ch_out[34]));
 sky130_fd_sc_hd__buf_6 wire51 (.A(net51),
    .X(ch_out[32]));
 sky130_fd_sc_hd__buf_6 wire52 (.A(net52),
    .X(ch_out[31]));
 sky130_fd_sc_hd__buf_6 wire53 (.A(net53),
    .X(ch_out[29]));
 sky130_fd_sc_hd__buf_6 wire54 (.A(net54),
    .X(ch_out[28]));
 sky130_fd_sc_hd__buf_6 wire55 (.A(net55),
    .X(ch_out[26]));
 sky130_fd_sc_hd__buf_6 wire56 (.A(net56),
    .X(ch_out[25]));
 sky130_fd_sc_hd__buf_6 wire57 (.A(net57),
    .X(ch_out[23]));
 sky130_fd_sc_hd__buf_6 wire58 (.A(net58),
    .X(ch_out[22]));
 sky130_fd_sc_hd__buf_6 wire59 (.A(net59),
    .X(ch_out[21]));
 sky130_fd_sc_hd__buf_4 wire6 (.A(net6),
    .X(ch_out[92]));
 sky130_fd_sc_hd__buf_6 wire60 (.A(net60),
    .X(ch_out[1]));
 sky130_fd_sc_hd__buf_6 wire61 (.A(net61),
    .X(ch_out[19]));
 sky130_fd_sc_hd__buf_6 wire62 (.A(net62),
    .X(ch_out[18]));
 sky130_fd_sc_hd__buf_6 wire63 (.A(net63),
    .X(ch_out[17]));
 sky130_fd_sc_hd__buf_6 wire64 (.A(net64),
    .X(ch_out[15]));
 sky130_fd_sc_hd__buf_6 wire65 (.A(net65),
    .X(ch_out[14]));
 sky130_fd_sc_hd__buf_6 wire66 (.A(net66),
    .X(ch_out[140]));
 sky130_fd_sc_hd__buf_6 wire67 (.A(net67),
    .X(ch_out[13]));
 sky130_fd_sc_hd__buf_6 wire68 (.A(net68),
    .X(ch_out[138]));
 sky130_fd_sc_hd__buf_6 wire69 (.A(net69),
    .X(ch_out[136]));
 sky130_fd_sc_hd__buf_4 wire7 (.A(net7),
    .X(ch_out[91]));
 sky130_fd_sc_hd__buf_6 wire70 (.A(net70),
    .X(ch_out[134]));
 sky130_fd_sc_hd__buf_6 wire71 (.A(net71),
    .X(ch_out[132]));
 sky130_fd_sc_hd__buf_6 wire72 (.A(net72),
    .X(ch_out[130]));
 sky130_fd_sc_hd__buf_6 wire73 (.A(net73),
    .X(ch_out[128]));
 sky130_fd_sc_hd__buf_6 wire74 (.A(net74),
    .X(ch_out[126]));
 sky130_fd_sc_hd__buf_6 wire75 (.A(net75),
    .X(ch_out[124]));
 sky130_fd_sc_hd__buf_6 wire76 (.A(net76),
    .X(ch_out[122]));
 sky130_fd_sc_hd__buf_6 wire77 (.A(net77),
    .X(ch_out[120]));
 sky130_fd_sc_hd__buf_6 wire78 (.A(net78),
    .X(ch_out[11]));
 sky130_fd_sc_hd__buf_6 wire79 (.A(net79),
    .X(ch_out[118]));
 sky130_fd_sc_hd__buf_4 wire8 (.A(net8),
    .X(ch_out[89]));
 sky130_fd_sc_hd__buf_6 wire80 (.A(net80),
    .X(ch_out[116]));
 sky130_fd_sc_hd__buf_6 wire81 (.A(net81),
    .X(ch_out[114]));
 sky130_fd_sc_hd__buf_6 wire82 (.A(net82),
    .X(ch_out[112]));
 sky130_fd_sc_hd__buf_6 wire83 (.A(net83),
    .X(ch_out[110]));
 sky130_fd_sc_hd__buf_6 wire84 (.A(net84),
    .X(ch_out[10]));
 sky130_fd_sc_hd__buf_6 wire85 (.A(net85),
    .X(ch_out[108]));
 sky130_fd_sc_hd__buf_6 wire86 (.A(net86),
    .X(ch_out[106]));
 sky130_fd_sc_hd__buf_4 wire87 (.A(net87),
    .X(ch_out[104]));
 sky130_fd_sc_hd__buf_4 wire88 (.A(net88),
    .X(ch_out[103]));
 sky130_fd_sc_hd__buf_4 wire89 (.A(net89),
    .X(ch_out[101]));
 sky130_fd_sc_hd__buf_4 wire9 (.A(net9),
    .X(ch_out[88]));
 sky130_fd_sc_hd__buf_4 wire90 (.A(net90),
    .X(ch_out[100]));
 sky130_fd_sc_hd__buf_6 wire91 (.A(net91),
    .X(ch_out[0]));
 sky130_fd_sc_hd__buf_4 wire92 (.A(ch_in[99]),
    .X(net92));
 sky130_fd_sc_hd__buf_4 wire93 (.A(ch_in[96]),
    .X(net93));
 sky130_fd_sc_hd__buf_4 wire94 (.A(ch_in[93]),
    .X(net94));
 sky130_fd_sc_hd__buf_4 wire95 (.A(ch_in[90]),
    .X(net95));
 sky130_fd_sc_hd__buf_6 wire96 (.A(ch_in[8]),
    .X(net96));
 sky130_fd_sc_hd__buf_4 wire97 (.A(ch_in[87]),
    .X(net97));
 sky130_fd_sc_hd__buf_4 wire98 (.A(ch_in[84]),
    .X(net98));
 sky130_fd_sc_hd__buf_4 wire99 (.A(ch_in[81]),
    .X(net99));
endmodule

