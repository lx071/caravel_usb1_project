VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO usb_top
  CLASS BLOCK ;
  FOREIGN usb_top ;
  ORIGIN 0.000 0.000 ;
  SIZE 500.000 BY 700.000 ;
  PIN app_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 308.760 4.000 309.360 ;
    END
  END app_clk
  PIN cfg_cska_usb[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 304.680 4.000 305.280 ;
    END
  END cfg_cska_usb[0]
  PIN cfg_cska_usb[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 303.320 4.000 303.920 ;
    END
  END cfg_cska_usb[1]
  PIN cfg_cska_usb[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END cfg_cska_usb[2]
  PIN cfg_cska_usb[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 300.600 4.000 301.200 ;
    END
  END cfg_cska_usb[3]
  PIN reg_ack
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 508.000 4.000 508.600 ;
    END
  END reg_ack
  PIN reg_addr[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.160 4.000 414.760 ;
    END
  END reg_addr[0]
  PIN reg_addr[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 412.800 4.000 413.400 ;
    END
  END reg_addr[1]
  PIN reg_addr[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END reg_addr[2]
  PIN reg_addr[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 410.080 4.000 410.680 ;
    END
  END reg_addr[3]
  PIN reg_addr[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 408.720 4.000 409.320 ;
    END
  END reg_addr[4]
  PIN reg_addr[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 407.360 4.000 407.960 ;
    END
  END reg_addr[5]
  PIN reg_addr[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 406.000 4.000 406.600 ;
    END
  END reg_addr[6]
  PIN reg_addr[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END reg_addr[7]
  PIN reg_addr[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 403.280 4.000 403.880 ;
    END
  END reg_addr[8]
  PIN reg_be[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 419.600 4.000 420.200 ;
    END
  END reg_be[0]
  PIN reg_be[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 418.240 4.000 418.840 ;
    END
  END reg_be[1]
  PIN reg_be[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.880 4.000 417.480 ;
    END
  END reg_be[2]
  PIN reg_be[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 415.520 4.000 416.120 ;
    END
  END reg_be[3]
  PIN reg_cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 400.560 4.000 401.160 ;
    END
  END reg_cs
  PIN reg_rdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END reg_rdata[0]
  PIN reg_rdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END reg_rdata[10]
  PIN reg_rdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 491.680 4.000 492.280 ;
    END
  END reg_rdata[11]
  PIN reg_rdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 490.320 4.000 490.920 ;
    END
  END reg_rdata[12]
  PIN reg_rdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 488.960 4.000 489.560 ;
    END
  END reg_rdata[13]
  PIN reg_rdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 487.600 4.000 488.200 ;
    END
  END reg_rdata[14]
  PIN reg_rdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END reg_rdata[15]
  PIN reg_rdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 484.880 4.000 485.480 ;
    END
  END reg_rdata[16]
  PIN reg_rdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 483.520 4.000 484.120 ;
    END
  END reg_rdata[17]
  PIN reg_rdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.160 4.000 482.760 ;
    END
  END reg_rdata[18]
  PIN reg_rdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 480.800 4.000 481.400 ;
    END
  END reg_rdata[19]
  PIN reg_rdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 505.280 4.000 505.880 ;
    END
  END reg_rdata[1]
  PIN reg_rdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 479.440 4.000 480.040 ;
    END
  END reg_rdata[20]
  PIN reg_rdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 478.080 4.000 478.680 ;
    END
  END reg_rdata[21]
  PIN reg_rdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.720 4.000 477.320 ;
    END
  END reg_rdata[22]
  PIN reg_rdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 475.360 4.000 475.960 ;
    END
  END reg_rdata[23]
  PIN reg_rdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 474.000 4.000 474.600 ;
    END
  END reg_rdata[24]
  PIN reg_rdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 472.640 4.000 473.240 ;
    END
  END reg_rdata[25]
  PIN reg_rdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 471.280 4.000 471.880 ;
    END
  END reg_rdata[26]
  PIN reg_rdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.920 4.000 470.520 ;
    END
  END reg_rdata[27]
  PIN reg_rdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 468.560 4.000 469.160 ;
    END
  END reg_rdata[28]
  PIN reg_rdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 467.200 4.000 467.800 ;
    END
  END reg_rdata[29]
  PIN reg_rdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 503.920 4.000 504.520 ;
    END
  END reg_rdata[2]
  PIN reg_rdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 465.840 4.000 466.440 ;
    END
  END reg_rdata[30]
  PIN reg_rdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 464.480 4.000 465.080 ;
    END
  END reg_rdata[31]
  PIN reg_rdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 502.560 4.000 503.160 ;
    END
  END reg_rdata[3]
  PIN reg_rdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 501.200 4.000 501.800 ;
    END
  END reg_rdata[4]
  PIN reg_rdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END reg_rdata[5]
  PIN reg_rdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 498.480 4.000 499.080 ;
    END
  END reg_rdata[6]
  PIN reg_rdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 497.120 4.000 497.720 ;
    END
  END reg_rdata[7]
  PIN reg_rdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 495.760 4.000 496.360 ;
    END
  END reg_rdata[8]
  PIN reg_rdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 494.400 4.000 495.000 ;
    END
  END reg_rdata[9]
  PIN reg_wdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 463.120 4.000 463.720 ;
    END
  END reg_wdata[0]
  PIN reg_wdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 449.520 4.000 450.120 ;
    END
  END reg_wdata[10]
  PIN reg_wdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 448.160 4.000 448.760 ;
    END
  END reg_wdata[11]
  PIN reg_wdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END reg_wdata[12]
  PIN reg_wdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END reg_wdata[13]
  PIN reg_wdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 444.080 4.000 444.680 ;
    END
  END reg_wdata[14]
  PIN reg_wdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 442.720 4.000 443.320 ;
    END
  END reg_wdata[15]
  PIN reg_wdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 441.360 4.000 441.960 ;
    END
  END reg_wdata[16]
  PIN reg_wdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 440.000 4.000 440.600 ;
    END
  END reg_wdata[17]
  PIN reg_wdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END reg_wdata[18]
  PIN reg_wdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 437.280 4.000 437.880 ;
    END
  END reg_wdata[19]
  PIN reg_wdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END reg_wdata[1]
  PIN reg_wdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.920 4.000 436.520 ;
    END
  END reg_wdata[20]
  PIN reg_wdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 434.560 4.000 435.160 ;
    END
  END reg_wdata[21]
  PIN reg_wdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 433.200 4.000 433.800 ;
    END
  END reg_wdata[22]
  PIN reg_wdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END reg_wdata[23]
  PIN reg_wdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 430.480 4.000 431.080 ;
    END
  END reg_wdata[24]
  PIN reg_wdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 429.120 4.000 429.720 ;
    END
  END reg_wdata[25]
  PIN reg_wdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 427.760 4.000 428.360 ;
    END
  END reg_wdata[26]
  PIN reg_wdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 426.400 4.000 427.000 ;
    END
  END reg_wdata[27]
  PIN reg_wdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 425.040 4.000 425.640 ;
    END
  END reg_wdata[28]
  PIN reg_wdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 423.680 4.000 424.280 ;
    END
  END reg_wdata[29]
  PIN reg_wdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 460.400 4.000 461.000 ;
    END
  END reg_wdata[2]
  PIN reg_wdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 422.320 4.000 422.920 ;
    END
  END reg_wdata[30]
  PIN reg_wdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 420.960 4.000 421.560 ;
    END
  END reg_wdata[31]
  PIN reg_wdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END reg_wdata[3]
  PIN reg_wdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 457.680 4.000 458.280 ;
    END
  END reg_wdata[4]
  PIN reg_wdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 456.320 4.000 456.920 ;
    END
  END reg_wdata[5]
  PIN reg_wdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 454.960 4.000 455.560 ;
    END
  END reg_wdata[6]
  PIN reg_wdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 453.600 4.000 454.200 ;
    END
  END reg_wdata[7]
  PIN reg_wdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END reg_wdata[8]
  PIN reg_wdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 450.880 4.000 451.480 ;
    END
  END reg_wdata[9]
  PIN reg_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.920 4.000 402.520 ;
    END
  END reg_wr
  PIN usb_clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 0.000 0.830 4.000 ;
    END
  END usb_clk
  PIN usb_in_dn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 696.000 1.750 700.000 ;
    END
  END usb_in_dn
  PIN usb_in_dp
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.550 696.000 0.830 700.000 ;
    END
  END usb_in_dp
  PIN usb_intr_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 5.150 696.000 5.430 700.000 ;
    END
  END usb_intr_o
  PIN usb_out_dn
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 696.000 3.590 700.000 ;
    END
  END usb_out_dn
  PIN usb_out_dp
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 696.000 2.670 700.000 ;
    END
  END usb_out_dp
  PIN usb_out_tx_oen
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 4.230 696.000 4.510 700.000 ;
    END
  END usb_out_tx_oen
  PIN usb_rstn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END usb_rstn
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 18.740 10.640 24.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 118.740 10.640 124.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 218.740 10.640 224.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 318.740 10.640 324.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 418.740 10.640 424.940 688.400 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 68.740 10.640 74.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 168.740 10.640 174.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 268.740 10.640 274.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 368.740 10.640 374.940 688.400 ;
    END
    PORT
      LAYER met4 ;
        RECT 468.740 10.640 474.940 688.400 ;
    END
  END vssd1
  PIN wbd_clk_int
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.040 4.000 306.640 ;
    END
  END wbd_clk_int
  PIN wbd_clk_usb
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 307.400 4.000 308.000 ;
    END
  END wbd_clk_usb
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 494.040 688.245 ;
      LAYER met1 ;
        RECT 0.530 4.460 494.040 690.840 ;
      LAYER met2 ;
        RECT 1.110 695.720 1.190 696.730 ;
        RECT 2.030 695.720 2.110 696.730 ;
        RECT 2.950 695.720 3.030 696.730 ;
        RECT 3.870 695.720 3.950 696.730 ;
        RECT 4.790 695.720 4.870 696.730 ;
        RECT 5.710 695.720 474.850 696.730 ;
        RECT 0.560 4.280 474.850 695.720 ;
        RECT 1.110 4.000 1.190 4.280 ;
        RECT 2.030 4.000 474.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 509.000 474.830 688.325 ;
        RECT 4.400 400.160 474.830 509.000 ;
        RECT 4.000 309.760 474.830 400.160 ;
        RECT 4.400 300.200 474.830 309.760 ;
        RECT 4.000 10.715 474.830 300.200 ;
      LAYER met4 ;
        RECT 9.495 137.535 18.340 669.625 ;
        RECT 25.340 137.535 68.340 669.625 ;
        RECT 75.340 137.535 118.340 669.625 ;
        RECT 125.340 137.535 168.340 669.625 ;
        RECT 175.340 137.535 218.340 669.625 ;
        RECT 225.340 137.535 268.340 669.625 ;
        RECT 275.340 137.535 318.340 669.625 ;
        RECT 325.340 137.535 329.985 669.625 ;
  END
END usb_top
END LIBRARY

